library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;

use work.cache_pack.all;

entity icache_tb is
end icache_tb;

architecture tb of icache_tb is

type adrs_buf_t is array (0 to 2047)  of std_logic_vector( 27 downto 0);

   signal rst   : std_logic;
   signal rst_46nsdel   : std_logic;
   signal clk125   : std_logic;
   signal clk200   : std_logic;

   signal a     : icache_i_t;
   signal y     : icache_o_t;
   signal ra    : icache_ram_o_t;
   signal ry    : icache_ram_i_t;
   signal ma    : mem_i_t;
   signal my    : mem_o_t;
   signal icccra : icccr_i_t;
   signal my_1delay : mem_o_t;
   signal ma_rdy_1wait_sig : std_logic;

   signal cavec  : std_logic_vector( 67 downto 0 );

   signal adrs_buf : adrs_buf_t;
   signal ack_pointer_thisc : std_logic_vector(10 downto 0);
   signal ack_pointer_thisr : std_logic_vector(10 downto 0);
   signal y_ack_1del_thisc : std_logic;
   signal y_ack_1del_thisr : std_logic;
begin

  --
  rst <= '1', '0' after 15 ns;
  rst_46nsdel <= rst after 46 ns;
  clk125 <= '0' after 4   ns when clk125 = '1' else '1' after 4   ns;
  clk200 <= '0' after 2.5 ns when clk200 = '1' else '1' after 2.5 ns;

-- .+....1....+....1....+....1....+....1....+....1....+....1....+....1....+....1
  dut : icache     port map ( rst => rst,
    clk125 => clk125, clk200 => clk200, a => a,
    y => y,           ra => ra,         ry => ry,
    ma => ma,         my => my ,        icccra => icccra );
  mem : configuration work.icache_ram_infer port map ( rst => rst,
    clk125 => clk125, 
    clk200 => clk200, ra => ry, ry => ra );

-- .+....1....+....1....+....1....+....1....+....1....+....1....+....1....+....1
  -- cache on/off selection
  -- --------------------------------------------------------------------------
    icccra.ic_onm <= '1'; -- cache on
--  icccra.ic_onm <= '0'; -- cache off
  -- --------------------------------------------------------------------------

  valid_rest : process( ack_pointer_thisr, y_ack_1del_thisr, rst_46nsdel)
  begin
    if(y_ack_1del_thisr = '1') and
      (ack_pointer_thisr(2 downto 0) = b"111") then
      a.a  <= x"aaaaaa0";
--    a.av <= '0';
      a.en <= '0';
    else
      a.a  <= adrs_buf(vtoi(ack_pointer_thisr));
--    a.av <= not rst_46nsdel;
      a.en <= not rst_46nsdel;
    end if;
  end process;

  ma.d <= (my.a(15 downto 2) & b"00" & my.a(15 downto 2) & b"10" ) and
   (
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack 
   ) ;

  my_1delay <= my after 5 ns;

  -- --------------------------------------------------------------------------
  gen_ready_1wait : process (my, my_1delay)
    variable mem_rdy_1wait : std_logic;
  begin
    if (my_1delay.en = '1') and
       (my.en        = '1') and
       (my_1delay.a = my.a) then mem_rdy_1wait := '1';
     else                        mem_rdy_1wait := '0';
     end if;
     ma_rdy_1wait_sig <=     mem_rdy_1wait;
  end process;
  -- --------------------------------------------------------------------------
  -- 1 wait
  ma.ack <= ma_rdy_1wait_sig;
  -- --------------------------------------------------------------------------

  ackfsm : process(ack_pointer_thisr, y.ack)
   variable ack_pointer_this : std_logic_vector(10 downto 0);
   variable y_ack_1del_this  : std_logic;
  begin
   ack_pointer_this := ack_pointer_thisr;
   y_ack_1del_this  := y_ack_1del_thisr;

   if(y.ack = '1') then
     ack_pointer_this := std_logic_vector(unsigned(ack_pointer_this) + 1);
   end if;
   y_ack_1del_this := y.ack;

   ack_pointer_thisc <= ack_pointer_this;
   y_ack_1del_thisc  <= y_ack_1del_this ;
  end process;

  p0_r0fsm : process(clk125, rst)
  begin
     if rst = '1' then
        ack_pointer_thisr <= b"000" & x"00";
        y_ack_1del_thisr  <= '0';
     elsif clk125 = '1' and clk125'event then
        ack_pointer_thisr <= ack_pointer_thisc;
        y_ack_1del_thisr  <= y_ack_1del_thisc ;
     end if;
  end process;


-- ---- access dump ------
  process
    file f0 : text is out "test.acc";
    variable l : line;
  begin

    wait for 1 ns;
    if(y.ack = '1') then
      hwrite(l, a.a );   write(l, string'(" "));
      hwrite(l, y.d );   write(l, string'(" "));
      -- write line --------------
      writeline(f0, l);
      deallocate(l);
    end if;
    wait for 7 ns;
  end process;

  -- test vector start
  -- read
  adrs_buf(   0) <= x"000010c";  -- miss
  adrs_buf(   1) <= x"000210a";  -- miss
  adrs_buf(   2) <= x"0004108";  -- miss
  adrs_buf(   3) <= x"0006106";  -- miss
  adrs_buf(   4) <= x"0001140";  -- miss
  adrs_buf(   5) <= x"0001158";
  adrs_buf(   6) <= x"0001176";  -- miss
  adrs_buf(   7) <= x"0201180";  -- miss
  adrs_buf(   8) <= x"03011a2";  -- miss
  adrs_buf(   9) <= x"04011c4";  -- miss
  adrs_buf(  10) <= x"05011e6";  -- miss
  adrs_buf(  11) <= x"000610e"; -- hit
  adrs_buf(  12) <= x"000115e"; -- hit
  adrs_buf(  13) <= x"000117e"; -- hit
  adrs_buf(  14) <= x"020119e"; -- hit
  adrs_buf(  15) <= x"03011be"; -- hit
  adrs_buf(  16) <= x"04011de"; -- hit
  adrs_buf(  17) <= x"05011fe"; -- hit
  adrs_buf(  18) <= x"0006100"; -- hit
  adrs_buf(  19) <= x"0001140"; -- hit
  adrs_buf(  20) <= x"0001160"; -- hit
  adrs_buf(  21) <= x"0201180"; -- hit
  adrs_buf(  22) <= x"03011a0"; -- hit
  adrs_buf(  23) <= x"04011c0"; -- hit
  adrs_buf(  24) <= x"05011e0"; -- hit
  adrs_buf(  25) <= x"021119e"; -- miss
  adrs_buf(  26) <= x"03111be"; -- miss
  adrs_buf(  27) <= x"04111de"; -- miss
  adrs_buf(  28) <= x"05111fe"; -- miss
  adrs_buf(  29) <= x"0000000";
  adrs_buf(  30) <= x"0000000";
  adrs_buf(  31) <= x"0000100"; -- miss
  adrs_buf(  32) <= x"000010e"; -- fill hit
  adrs_buf(  33) <= x"0000000";
  adrs_buf(  34) <= x"0002100"; -- miss
  adrs_buf(  35) <= x"000210c"; -- fill hit
  adrs_buf(  36) <= x"0000000";
  adrs_buf(  37) <= x"0000100"; -- miss
  adrs_buf(  38) <= x"000010a"; -- fill hit
  adrs_buf(  39) <= x"0000000";
  adrs_buf(  40) <= x"0002100"; -- miss
  adrs_buf(  41) <= x"0002108"; -- fill hit
  adrs_buf(  42) <= x"0000000";
  adrs_buf(  43) <= x"0000100"; -- miss
  adrs_buf(  44) <= x"0000106"; -- fill hit
  adrs_buf(  45) <= x"0000000";
  adrs_buf(  46) <= x"0002100"; -- miss
  adrs_buf(  47) <= x"0002104"; -- fill hit
  adrs_buf(  48) <= x"0000000";
  adrs_buf(  49) <= x"0000100"; -- miss
  adrs_buf(  50) <= x"0000102"; -- fill hit
  adrs_buf(  51) <= x"0000000";
  adrs_buf(  52) <= x"0002100"; -- miss 
  adrs_buf(  53) <= x"0002100"; -- fill hit
  adrs_buf(  54) <= x"0000000";
  adrs_buf(  55) <= x"000820e"; -- miss
  adrs_buf(  56) <= x"0008200"; -- fill hit
  adrs_buf(  57) <= x"0000000";
  adrs_buf(  58) <= x"000420e"; -- miss
  adrs_buf(  59) <= x"0004204"; -- fill hit
  adrs_buf(  60) <= x"0000000";
  adrs_buf(  61) <= x"000820e"; -- miss
  adrs_buf(  62) <= x"0008208"; -- fill hit
  adrs_buf(  63) <= x"0000000";
  adrs_buf(  64) <= x"000420e"; -- miss
  adrs_buf(  65) <= x"000420c"; -- fill hit
  adrs_buf(  66) <= x"0000000";
  adrs_buf(  67) <= x"000820e"; -- miss
  adrs_buf(  68) <= x"0008210"; -- fill hit
  adrs_buf(  69) <= x"0000000";
  adrs_buf(  70) <= x"000420e"; -- miss
  adrs_buf(  71) <= x"0004214"; -- fill hit
  adrs_buf(  72) <= x"0000000";
  adrs_buf(  73) <= x"000820e"; -- miss
  adrs_buf(  74) <= x"0008218"; -- fill hit
  adrs_buf(  75) <= x"0000000";
  adrs_buf(  76) <= x"000420e"; -- miss
  adrs_buf(  77) <= x"000421c"; -- fill hit
  adrs_buf(  78) <= x"0000000";
  adrs_buf(  79) <= x"000820e"; -- miss
  adrs_buf(  80) <= x"000820e"; -- fill hit
  adrs_buf(  81) <= x"0000000";
  adrs_buf(  82) <= x"ffffff0"; -- miss
  adrs_buf(  83) <= x"0000000";
  adrs_buf(  84) <= x"0004200"; -- miss
  adrs_buf(  85) <= x"0004204"; -- fill hit no wait
  adrs_buf(  86) <= x"000421e"; -- fill hit wait
  adrs_buf(  87) <= x"0000000";
  adrs_buf(  88) <= x"0008200"; -- miss
  adrs_buf(  89) <= x"0008202"; -- fill hit no wait
  adrs_buf(  90) <= x"000821c"; -- fill hit wait
  adrs_buf(  91) <= x"0000000";
  adrs_buf(  92) <= x"0004218"; -- miss
  adrs_buf(  93) <= x"000421c"; -- fill hit no wait
  adrs_buf(  94) <= x"0004216"; -- fill hit wait
  adrs_buf(  95) <= x"0000000";
  adrs_buf(  96) <= x"0000206"; -- corner case 4n+2 same
  adrs_buf(  97) <= x"0000206";
  adrs_buf(  98) <= x"0000206";
  adrs_buf(  99) <= x"0000206";
  adrs_buf( 100) <= x"0000206";
  adrs_buf( 101) <= x"0000210";
  adrs_buf( 102) <= x"0000210";
  adrs_buf( 103) <= x"0000210";
  adrs_buf( 104) <= x"0000210";
  adrs_buf( 105) <= x"0000210";
  adrs_buf( 106) <= x"0000212";
  adrs_buf( 107) <= x"0000212";
  adrs_buf( 108) <= x"0000212";
  adrs_buf( 109) <= x"0000212";
  adrs_buf( 110) <= x"0000212";
  adrs_buf( 111) <= x"0000000";
  adrs_buf( 112) <= x"0000000";
  adrs_buf( 113) <= x"0000000";
  adrs_buf( 114) <= x"0000000";
  adrs_buf( 115) <= x"0000000";
  adrs_buf( 116) <= x"0000000";
  adrs_buf( 117) <= x"0000000";
  adrs_buf( 118) <= x"0000000";
  adrs_buf( 119) <= x"0000000";
  adrs_buf( 120) <= x"0000000";
  adrs_buf( 121) <= x"0000000";
  adrs_buf( 122) <= x"0000000";
  adrs_buf( 123) <= x"0000000";
  adrs_buf( 124) <= x"0000000";
  adrs_buf( 125) <= x"0000000";
  adrs_buf( 126) <= x"00013e0";
  adrs_buf( 127) <= x"00013e2";
  adrs_buf( 128) <= x"00013e4";
  adrs_buf( 129) <= x"00013e6";
  adrs_buf( 130) <= x"00013e8";
  adrs_buf( 131) <= x"00013ea";
  adrs_buf( 132) <= x"00013ec";
  adrs_buf( 133) <= x"00013ee";
  adrs_buf( 134) <= x"00013f0";
  adrs_buf( 135) <= x"00013f2";
  adrs_buf( 136) <= x"00013f4";
  adrs_buf( 137) <= x"00013f6";
  adrs_buf( 138) <= x"00013f8";
  adrs_buf( 139) <= x"00013fe";
  adrs_buf( 140) <= x"0001400";
  adrs_buf( 141) <= x"0001402";
  adrs_buf( 142) <= x"0001404";
  adrs_buf( 143) <= x"0001406";
  adrs_buf( 144) <= x"0001408";
  adrs_buf( 145) <= x"000140a";
  adrs_buf( 146) <= x"000140c";
  adrs_buf( 147) <= x"000140e";
  adrs_buf( 148) <= x"0001410";
  adrs_buf( 149) <= x"0001416";
  adrs_buf( 150) <= x"0001418";
  adrs_buf( 151) <= x"000141a";
  adrs_buf( 152) <= x"000141c";
  adrs_buf( 153) <= x"000141e";
  adrs_buf( 154) <= x"0001420";
  adrs_buf( 155) <= x"0001422";
  adrs_buf( 156) <= x"0001424";
  adrs_buf( 157) <= x"0001426";
  adrs_buf( 158) <= x"000143c";
  adrs_buf( 159) <= x"000143e";
  adrs_buf( 160) <= x"0001440";
  adrs_buf( 161) <= x"0001442";
  adrs_buf( 162) <= x"0001428";
  adrs_buf( 163) <= x"000142a";
  adrs_buf( 164) <= x"000142c";
  adrs_buf( 165) <= x"000142e";
  adrs_buf( 166) <= x"0001430";
  adrs_buf( 167) <= x"0001432";
  adrs_buf( 168) <= x"0001434";
  adrs_buf( 169) <= x"0001436";
  adrs_buf( 170) <= x"0001438";
  adrs_buf( 171) <= x"000143a";
  adrs_buf( 172) <= x"0001444";
  adrs_buf( 173) <= x"0001446";
  adrs_buf( 174) <= x"0001448";
  adrs_buf( 175) <= x"000144a";
  adrs_buf( 176) <= x"000144c";
  adrs_buf( 177) <= x"000145e";
  adrs_buf( 178) <= x"0001460";
  adrs_buf( 179) <= x"0001462";
  adrs_buf( 180) <= x"0001464";
  adrs_buf( 181) <= x"0001466";
  adrs_buf( 182) <= x"0001468";
  adrs_buf( 183) <= x"000146a";
  adrs_buf( 184) <= x"0001478";
  adrs_buf( 185) <= x"000147a";
  adrs_buf( 186) <= x"000147c";
  adrs_buf( 187) <= x"000147e";
  adrs_buf( 188) <= x"0001486";
  adrs_buf( 189) <= x"0001488";
  adrs_buf( 190) <= x"000148a";
  adrs_buf( 191) <= x"000148c";
  adrs_buf( 192) <= x"000148e";
  adrs_buf( 193) <= x"0001490";
  adrs_buf( 194) <= x"0001480";
  adrs_buf( 195) <= x"0001482";
  adrs_buf( 196) <= x"0001484";
  adrs_buf( 197) <= x"000146c";
  adrs_buf( 198) <= x"000146e";
  adrs_buf( 199) <= x"0001470";
  adrs_buf( 200) <= x"0001472";
  adrs_buf( 201) <= x"0001474";
  adrs_buf( 202) <= x"0001476";
  adrs_buf( 203) <= x"0001492";
  adrs_buf( 204) <= x"0001494";
  adrs_buf( 205) <= x"0001496";
  adrs_buf( 206) <= x"0001498";
  adrs_buf( 207) <= x"000149a";
  adrs_buf( 208) <= x"000149c";
  adrs_buf( 209) <= x"000149e";
  adrs_buf( 210) <= x"00014a0";
  adrs_buf( 211) <= x"00014a2";
  adrs_buf( 212) <= x"00014a4";
  adrs_buf( 213) <= x"00014a6";
  adrs_buf( 214) <= x"00014a8";
  adrs_buf( 215) <= x"00014aa";
  adrs_buf( 216) <= x"00014ac";
  adrs_buf( 217) <= x"00014ae";
  adrs_buf( 218) <= x"00014b0";
  adrs_buf( 219) <= x"00014b2";
  adrs_buf( 220) <= x"00014b4";
  adrs_buf( 221) <= x"00014b6";
  adrs_buf( 222) <= x"00014b8";
  adrs_buf( 223) <= x"00014ba";
  adrs_buf( 224) <= x"00014bc";
  adrs_buf( 225) <= x"00014be";
  adrs_buf( 226) <= x"00014c0";
  adrs_buf( 227) <= x"00014c2";
  adrs_buf( 228) <= x"00014c4";
  adrs_buf( 229) <= x"00014c6";
  adrs_buf( 230) <= x"00014c8";
  adrs_buf( 231) <= x"00014ca";
  adrs_buf( 232) <= x"00014cc";
  adrs_buf( 233) <= x"00014ce";
  adrs_buf( 234) <= x"00014d0";
  adrs_buf( 235) <= x"00014d2";
  adrs_buf( 236) <= x"00014d4";
  adrs_buf( 237) <= x"00014d6";
  adrs_buf( 238) <= x"00014d8";
  adrs_buf( 239) <= x"00014da";
  adrs_buf( 240) <= x"00014dc";
  adrs_buf( 241) <= x"00014de";
  adrs_buf( 242) <= x"00014e0";
  adrs_buf( 243) <= x"00014e2";
  adrs_buf( 244) <= x"00014e4";
  adrs_buf( 245) <= x"00014e6";
  adrs_buf( 246) <= x"00014e8";
  adrs_buf( 247) <= x"00014ea";
  adrs_buf( 248) <= x"00014ec";
  adrs_buf( 249) <= x"00014ee";
  adrs_buf( 250) <= x"00014f0";
  adrs_buf( 251) <= x"00014f2";
  adrs_buf( 252) <= x"00014f4";
  adrs_buf( 253) <= x"00014f6";
  adrs_buf( 254) <= x"00014f8";
  adrs_buf( 255) <= x"00014fa";
  adrs_buf( 256) <= x"00014fc";
  adrs_buf( 257) <= x"00014fe";
  adrs_buf( 258) <= x"0001500";
  adrs_buf( 259) <= x"0001502";
  adrs_buf( 260) <= x"0001504";
  adrs_buf( 261) <= x"0001506";
  adrs_buf( 262) <= x"0001508";
  adrs_buf( 263) <= x"000150a";
  adrs_buf( 264) <= x"000150c";
  adrs_buf( 265) <= x"000150e";
  adrs_buf( 266) <= x"0001510";
  adrs_buf( 267) <= x"0001512";
  adrs_buf( 268) <= x"0001514";
  adrs_buf( 269) <= x"0001516";
  adrs_buf( 270) <= x"0001518";
  adrs_buf( 271) <= x"000151a";
  adrs_buf( 272) <= x"000151c";
  adrs_buf( 273) <= x"000151e";
  adrs_buf( 274) <= x"0001520";
  adrs_buf( 275) <= x"0001522";
  adrs_buf( 276) <= x"0001524";
  adrs_buf( 277) <= x"0001526";
  adrs_buf( 278) <= x"0001528";
  adrs_buf( 279) <= x"000152a";
  adrs_buf( 280) <= x"000152c";
  adrs_buf( 281) <= x"000152e";
  adrs_buf( 282) <= x"0001530";
  adrs_buf( 283) <= x"0001532";
  adrs_buf( 284) <= x"0001534";
  adrs_buf( 285) <= x"0001536";
  adrs_buf( 286) <= x"0001538";
  adrs_buf( 287) <= x"000153a";
  adrs_buf( 288) <= x"000153c";
  adrs_buf( 289) <= x"000153e";
  adrs_buf( 290) <= x"0001544";
  adrs_buf( 291) <= x"0001546";
  adrs_buf( 292) <= x"000156c";
  adrs_buf( 293) <= x"000156e";
  adrs_buf( 294) <= x"0001570";
  adrs_buf( 295) <= x"0001572";
  adrs_buf( 296) <= x"0001574";
  adrs_buf( 297) <= x"0001576";
  adrs_buf( 298) <= x"0000126";
  adrs_buf( 299) <= x"0000128";
  adrs_buf( 300) <= x"000012a";
  adrs_buf( 301) <= x"00015a0";
  adrs_buf( 302) <= x"00015a2";
  adrs_buf( 303) <= x"00015a4";
  adrs_buf( 304) <= x"00015a6";
  adrs_buf( 305) <= x"00015ac";
  adrs_buf( 306) <= x"00015ae";
  adrs_buf( 307) <= x"00015b0";
  adrs_buf( 308) <= x"00015b2";
  adrs_buf( 309) <= x"00015b4";
  adrs_buf( 310) <= x"00015b6";
  adrs_buf( 311) <= x"00015b8";
  adrs_buf( 312) <= x"00015ba";
  adrs_buf( 313) <= x"00015bc";
  adrs_buf( 314) <= x"00015be";
  adrs_buf( 315) <= x"00015c0";
  adrs_buf( 316) <= x"00015c2";
  adrs_buf( 317) <= x"00015c4";
  adrs_buf( 318) <= x"00015c6";
  adrs_buf( 319) <= x"00015c8";
  adrs_buf( 320) <= x"00015ca";
  adrs_buf( 321) <= x"00015cc";
  adrs_buf( 322) <= x"00015ce";
  adrs_buf( 323) <= x"00015d0";
  adrs_buf( 324) <= x"00015d2";
  adrs_buf( 325) <= x"00015d4";
  adrs_buf( 326) <= x"00015d6";
  adrs_buf( 327) <= x"00015d8";
  adrs_buf( 328) <= x"00015da";
  adrs_buf( 329) <= x"00015dc";
  adrs_buf( 330) <= x"00015de";
  adrs_buf( 331) <= x"00015e0";
  adrs_buf( 332) <= x"00015e2";
  adrs_buf( 333) <= x"00015e4";
  adrs_buf( 334) <= x"00015e6";
  adrs_buf( 335) <= x"00015e8";
  adrs_buf( 336) <= x"00015ea";
  adrs_buf( 337) <= x"00015ec";
  adrs_buf( 338) <= x"00015ee";
  adrs_buf( 339) <= x"00015f0";
  adrs_buf( 340) <= x"00015f2";
  adrs_buf( 341) <= x"00015f4";
  adrs_buf( 342) <= x"00015f6";
  adrs_buf( 343) <= x"00015f8";
  adrs_buf( 344) <= x"00015fa";
  adrs_buf( 345) <= x"00015fc";
  adrs_buf( 346) <= x"00015fe";
  adrs_buf( 347) <= x"0001600";
  adrs_buf( 348) <= x"0001602";
  adrs_buf( 349) <= x"0001604";
  adrs_buf( 350) <= x"0001606";
  adrs_buf( 351) <= x"0001608";
  adrs_buf( 352) <= x"000160a";
  adrs_buf( 353) <= x"000160c";
  adrs_buf( 354) <= x"000160e";
  adrs_buf( 355) <= x"0001610";
  adrs_buf( 356) <= x"0001612";
  adrs_buf( 357) <= x"0001614";
  adrs_buf( 358) <= x"0001616";
  adrs_buf( 359) <= x"0001618";
  adrs_buf( 360) <= x"000161a";
  adrs_buf( 361) <= x"000161c";
  adrs_buf( 362) <= x"000161e";
  adrs_buf( 363) <= x"0001620";
  adrs_buf( 364) <= x"0001622";
  adrs_buf( 365) <= x"0001624";
  adrs_buf( 366) <= x"0001626";
  adrs_buf( 367) <= x"0001628";
  adrs_buf( 368) <= x"000162a";
  adrs_buf( 369) <= x"000162c";
  adrs_buf( 370) <= x"000162e";
  adrs_buf( 371) <= x"0001630";
  adrs_buf( 372) <= x"0001632";
  adrs_buf( 373) <= x"0001634";
  adrs_buf( 374) <= x"0001636";
  adrs_buf( 375) <= x"0001638";
  adrs_buf( 376) <= x"000163a";
  adrs_buf( 377) <= x"000163c";
  adrs_buf( 378) <= x"000163e";
  adrs_buf( 379) <= x"0001640";
  adrs_buf( 380) <= x"0001642";
  adrs_buf( 381) <= x"0001644";
  adrs_buf( 382) <= x"0001646";
  adrs_buf( 383) <= x"0001648";
  adrs_buf( 384) <= x"000164a";
  adrs_buf( 385) <= x"000164c";
  adrs_buf( 386) <= x"000164e";
  adrs_buf( 387) <= x"0001650";
  adrs_buf( 388) <= x"0001652";
  adrs_buf( 389) <= x"0001654";
  adrs_buf( 390) <= x"0001656";
  adrs_buf( 391) <= x"0001658";
  adrs_buf( 392) <= x"000165a";
  adrs_buf( 393) <= x"000165c";
  adrs_buf( 394) <= x"000165e";
  adrs_buf( 395) <= x"0001660";
  adrs_buf( 396) <= x"0001662";
  adrs_buf( 397) <= x"0001664";
  adrs_buf( 398) <= x"0001666";
  adrs_buf( 399) <= x"0001668";
  adrs_buf( 400) <= x"000166a";
  adrs_buf( 401) <= x"000166c";
  adrs_buf( 402) <= x"000166e";
  adrs_buf( 403) <= x"0001670";
  adrs_buf( 404) <= x"0001672";
  adrs_buf( 405) <= x"0001674";
  adrs_buf( 406) <= x"0001676";
  adrs_buf( 407) <= x"0001678";
  adrs_buf( 408) <= x"000167a";
  adrs_buf( 409) <= x"000167c";
  adrs_buf( 410) <= x"000167e";
  adrs_buf( 411) <= x"0001680";
  adrs_buf( 412) <= x"0001682";
  adrs_buf( 413) <= x"0001684";
  adrs_buf( 414) <= x"0001686";
  adrs_buf( 415) <= x"0001688";
  adrs_buf( 416) <= x"000168a";
  adrs_buf( 417) <= x"000168c";
  adrs_buf( 418) <= x"000168e";
  adrs_buf( 419) <= x"0001690";
  adrs_buf( 420) <= x"0001692";
  adrs_buf( 421) <= x"0001694";
  adrs_buf( 422) <= x"0001696";
  adrs_buf( 423) <= x"0001698";
  adrs_buf( 424) <= x"000169a";
  adrs_buf( 425) <= x"000169c";
  adrs_buf( 426) <= x"000169e";
  adrs_buf( 427) <= x"00016a0";
  adrs_buf( 428) <= x"00016a2";
  adrs_buf( 429) <= x"00016a4";
  adrs_buf( 430) <= x"00016a6";
  adrs_buf( 431) <= x"00016a8";
  adrs_buf( 432) <= x"00016aa";
  adrs_buf( 433) <= x"00016ac";
  adrs_buf( 434) <= x"00016ae";
  adrs_buf( 435) <= x"00016b0";
  adrs_buf( 436) <= x"00016b2";
  adrs_buf( 437) <= x"00016b4";
  adrs_buf( 438) <= x"00016b6";
  adrs_buf( 439) <= x"00016b8";
  adrs_buf( 440) <= x"00016ba";
  adrs_buf( 441) <= x"00016bc";
  adrs_buf( 442) <= x"00016be";
  adrs_buf( 443) <= x"00016c0";
  adrs_buf( 444) <= x"00016c2";
  adrs_buf( 445) <= x"00016c4";
  adrs_buf( 446) <= x"00016c6";
  adrs_buf( 447) <= x"00016c8";
  adrs_buf( 448) <= x"00016ca";
  adrs_buf( 449) <= x"00016cc";
  adrs_buf( 450) <= x"00016ce";
  adrs_buf( 451) <= x"00016d0";
  adrs_buf( 452) <= x"00016d2";
  adrs_buf( 453) <= x"00016d4";
  adrs_buf( 454) <= x"00016d6";
  adrs_buf( 455) <= x"00016d8";
  adrs_buf( 456) <= x"00016da";
  adrs_buf( 457) <= x"00016dc";
  adrs_buf( 458) <= x"00016de";
  adrs_buf( 459) <= x"00016e0";
  adrs_buf( 460) <= x"00016e2";
  adrs_buf( 461) <= x"00016e4";
  adrs_buf( 462) <= x"00016e6";
  adrs_buf( 463) <= x"00016e8";
  adrs_buf( 464) <= x"00016ea";
  adrs_buf( 465) <= x"00016ec";
  adrs_buf( 466) <= x"00016ee";
  adrs_buf( 467) <= x"00016f0";
  adrs_buf( 468) <= x"00016f2";
  adrs_buf( 469) <= x"00016f4";
  adrs_buf( 470) <= x"00016f6";
  adrs_buf( 471) <= x"00016f8";
  adrs_buf( 472) <= x"00016fa";
  adrs_buf( 473) <= x"00016fc";
  adrs_buf( 474) <= x"00016fe";
  adrs_buf( 475) <= x"0001700";
  adrs_buf( 476) <= x"0001702";
  adrs_buf( 477) <= x"0001704";
  adrs_buf( 478) <= x"0001706";
  adrs_buf( 479) <= x"0001708";
  adrs_buf( 480) <= x"000170a";
  adrs_buf( 481) <= x"000170c";
  adrs_buf( 482) <= x"000170e";
  adrs_buf( 483) <= x"0001710";
  adrs_buf( 484) <= x"0001712";
  adrs_buf( 485) <= x"0001714";
  adrs_buf( 486) <= x"0001716";
  adrs_buf( 487) <= x"0001718";
  adrs_buf( 488) <= x"000171a";
  adrs_buf( 489) <= x"000171c";
  adrs_buf( 490) <= x"000171e";
  adrs_buf( 491) <= x"0001720";
  adrs_buf( 492) <= x"0001722";
  adrs_buf( 493) <= x"0001724";
  adrs_buf( 494) <= x"0001726";
  adrs_buf( 495) <= x"0001728";
  adrs_buf( 496) <= x"000172a";
  adrs_buf( 497) <= x"000172c";
  adrs_buf( 498) <= x"000172e";
  adrs_buf( 499) <= x"0001730";
  adrs_buf( 500) <= x"0001732";
  adrs_buf( 501) <= x"0001734";
  adrs_buf( 502) <= x"0001736";
  adrs_buf( 503) <= x"0001738";
  adrs_buf( 504) <= x"000173a";
  adrs_buf( 505) <= x"000173c";
  adrs_buf( 506) <= x"000173e";
  adrs_buf( 507) <= x"0001740";
  adrs_buf( 508) <= x"0001742";
  adrs_buf( 509) <= x"0001744";
  adrs_buf( 510) <= x"0001746";
  adrs_buf( 511) <= x"0001748";
  adrs_buf( 512) <= x"000174a";
  adrs_buf( 513) <= x"000174c";
  adrs_buf( 514) <= x"000174e";
  adrs_buf( 515) <= x"0001750";
  adrs_buf( 516) <= x"0001752";
  adrs_buf( 517) <= x"0001754";
  adrs_buf( 518) <= x"0001756";
  adrs_buf( 519) <= x"0001758";
  adrs_buf( 520) <= x"000175a";
  adrs_buf( 521) <= x"000175c";
  adrs_buf( 522) <= x"000175e";
  adrs_buf( 523) <= x"0001760";
  adrs_buf( 524) <= x"0001762";
  adrs_buf( 525) <= x"0001764";
  adrs_buf( 526) <= x"0001766";
  adrs_buf( 527) <= x"0001768";
  adrs_buf( 528) <= x"000176a";
  adrs_buf( 529) <= x"000176c";
  adrs_buf( 530) <= x"000176e";
  adrs_buf( 531) <= x"0001770";
  adrs_buf( 532) <= x"0001772";
  adrs_buf( 533) <= x"0001774";
  adrs_buf( 534) <= x"0001776";
  adrs_buf( 535) <= x"0001778";
  adrs_buf( 536) <= x"000177a";
  adrs_buf( 537) <= x"000177c";
  adrs_buf( 538) <= x"000177e";
  adrs_buf( 539) <= x"0001780";
  adrs_buf( 540) <= x"0001782";
  adrs_buf( 541) <= x"0001784";
  adrs_buf( 542) <= x"0001786";
  adrs_buf( 543) <= x"0001788";
  adrs_buf( 544) <= x"000178a";
  adrs_buf( 545) <= x"000178c";
  adrs_buf( 546) <= x"000178e";
  adrs_buf( 547) <= x"0001790";
  adrs_buf( 548) <= x"0001792";
  adrs_buf( 549) <= x"0001794";
  adrs_buf( 550) <= x"0001796";
  adrs_buf( 551) <= x"0001798";
  adrs_buf( 552) <= x"000179a";
  adrs_buf( 553) <= x"000179c";
  adrs_buf( 554) <= x"000179e";
  adrs_buf( 555) <= x"00017a0";
  adrs_buf( 556) <= x"00017a2";
  adrs_buf( 557) <= x"00017a4";
  adrs_buf( 558) <= x"00017a6";
  adrs_buf( 559) <= x"00017a8";
  adrs_buf( 560) <= x"00017aa";
  adrs_buf( 561) <= x"00017ac";
  adrs_buf( 562) <= x"00017ae";
  adrs_buf( 563) <= x"00017b0";
  adrs_buf( 564) <= x"00017b2";
  adrs_buf( 565) <= x"00017b4";
  adrs_buf( 566) <= x"00017b6";
  adrs_buf( 567) <= x"00017b8";
  adrs_buf( 568) <= x"00017ba";
  adrs_buf( 569) <= x"00017bc";
  adrs_buf( 570) <= x"00017be";
  adrs_buf( 571) <= x"00017c0";
  adrs_buf( 572) <= x"00017c2";
  adrs_buf( 573) <= x"00017c4";
  adrs_buf( 574) <= x"00017c6";
  adrs_buf( 575) <= x"00017c8";
  adrs_buf( 576) <= x"00017ca";
  adrs_buf( 577) <= x"00017cc";
  adrs_buf( 578) <= x"00017ce";
  adrs_buf( 579) <= x"00017d0";
  adrs_buf( 580) <= x"00017d2";
  adrs_buf( 581) <= x"00017d4";
  adrs_buf( 582) <= x"00017d6";
  adrs_buf( 583) <= x"00017d8";
  adrs_buf( 584) <= x"00017da";
  adrs_buf( 585) <= x"00017dc";
  adrs_buf( 586) <= x"00017de";
  adrs_buf( 587) <= x"00017e0";
  adrs_buf( 588) <= x"00017e2";
  adrs_buf( 589) <= x"00017e4";
  adrs_buf( 590) <= x"00017e6";
  adrs_buf( 591) <= x"00017e8";
  adrs_buf( 592) <= x"00017ea";
  adrs_buf( 593) <= x"00017ec";
  adrs_buf( 594) <= x"00017ee";
  adrs_buf( 595) <= x"00017f0";
  adrs_buf( 596) <= x"00017f2";
  adrs_buf( 597) <= x"00017f4";
  adrs_buf( 598) <= x"00017f6";
  adrs_buf( 599) <= x"00017f8";
  adrs_buf( 600) <= x"00017fa";
  adrs_buf( 601) <= x"00017fc";
  adrs_buf( 602) <= x"00017fe";
  adrs_buf( 603) <= x"0001800";
  adrs_buf( 604) <= x"0001802";
  adrs_buf( 605) <= x"0001804";
  adrs_buf( 606) <= x"0001806";
  adrs_buf( 607) <= x"0001808";
  adrs_buf( 608) <= x"000180a";
  adrs_buf( 609) <= x"000180c";
  adrs_buf( 610) <= x"000180e";
  adrs_buf( 611) <= x"0001810";
  adrs_buf( 612) <= x"0001812";
  adrs_buf( 613) <= x"0001814";
  adrs_buf( 614) <= x"0001816";
  adrs_buf( 615) <= x"0001818";
  adrs_buf( 616) <= x"000181a";
  adrs_buf( 617) <= x"000181c";
  adrs_buf( 618) <= x"000181e";
  adrs_buf( 619) <= x"0001820";
  adrs_buf( 620) <= x"0001822";
  adrs_buf( 621) <= x"0001824";
  adrs_buf( 622) <= x"0001826";
  adrs_buf( 623) <= x"0001828";
  adrs_buf( 624) <= x"000182a";
  adrs_buf( 625) <= x"000182c";
  adrs_buf( 626) <= x"000182e";
  adrs_buf( 627) <= x"0001830";
  adrs_buf( 628) <= x"0001832";
  adrs_buf( 629) <= x"0001834";
  adrs_buf( 630) <= x"0001836";
  adrs_buf( 631) <= x"0001838";
  adrs_buf( 632) <= x"000183a";
  adrs_buf( 633) <= x"000183c";
  adrs_buf( 634) <= x"000183e";
  adrs_buf( 635) <= x"0001840";
  adrs_buf( 636) <= x"0001842";
  adrs_buf( 637) <= x"0001844";
  adrs_buf( 638) <= x"0001846";
  adrs_buf( 639) <= x"0001848";
  adrs_buf( 640) <= x"000184a";
  adrs_buf( 641) <= x"000184c";
  adrs_buf( 642) <= x"000184e";
  adrs_buf( 643) <= x"0001850";
  adrs_buf( 644) <= x"0001852";
  adrs_buf( 645) <= x"0001854";
  adrs_buf( 646) <= x"0001856";
  adrs_buf( 647) <= x"0001858";
  adrs_buf( 648) <= x"000185a";
  adrs_buf( 649) <= x"000185c";
  adrs_buf( 650) <= x"000185e";
  adrs_buf( 651) <= x"0001860";
  adrs_buf( 652) <= x"0001862";
  adrs_buf( 653) <= x"0001864";
  adrs_buf( 654) <= x"0001866";
  adrs_buf( 655) <= x"0001868";
  adrs_buf( 656) <= x"000186a";
  adrs_buf( 657) <= x"000186c";
  adrs_buf( 658) <= x"000186e";
  adrs_buf( 659) <= x"0001870";
  adrs_buf( 660) <= x"0001872";
  adrs_buf( 661) <= x"0001874";
  adrs_buf( 662) <= x"0001876";
  adrs_buf( 663) <= x"0001878";
  adrs_buf( 664) <= x"000187a";
  adrs_buf( 665) <= x"000187c";
  adrs_buf( 666) <= x"000187e";
  adrs_buf( 667) <= x"0001880";
  adrs_buf( 668) <= x"0001882";
  adrs_buf( 669) <= x"0001884";
  adrs_buf( 670) <= x"0001886";
  adrs_buf( 671) <= x"0001888";
  adrs_buf( 672) <= x"000188a";
  adrs_buf( 673) <= x"00018d8";
  adrs_buf( 674) <= x"00018da";
  adrs_buf( 675) <= x"00018dc";
  adrs_buf( 676) <= x"00018de";
  adrs_buf( 677) <= x"00018e0";
  adrs_buf( 678) <= x"00018e2";
  adrs_buf( 679) <= x"000012c";
  adrs_buf( 680) <= x"000012e";
  adrs_buf( 681) <= x"0000130";
  adrs_buf( 682) <= x"0001910";
  adrs_buf( 683) <= x"0001912";
  adrs_buf( 684) <= x"0001914";
  adrs_buf( 685) <= x"0001916";
  adrs_buf( 686) <= x"000191c";
  adrs_buf( 687) <= x"000191e";
  adrs_buf( 688) <= x"0001920";
  adrs_buf( 689) <= x"0001922";
  adrs_buf( 690) <= x"0001930";
  adrs_buf( 691) <= x"0001932";
  adrs_buf( 692) <= x"0001938";
  adrs_buf( 693) <= x"000193a";
  adrs_buf( 694) <= x"0001940";
  adrs_buf( 695) <= x"0001942";
  adrs_buf( 696) <= x"0001944";
  adrs_buf( 697) <= x"0001946";
  adrs_buf( 698) <= x"0001948";
  adrs_buf( 699) <= x"000194a";
  adrs_buf( 700) <= x"000194c";
  adrs_buf( 701) <= x"000194e";
  adrs_buf( 702) <= x"0001950";
  adrs_buf( 703) <= x"0001952";
  adrs_buf( 704) <= x"0001954";
  adrs_buf( 705) <= x"0001956";
  adrs_buf( 706) <= x"0001958";
  adrs_buf( 707) <= x"000195a";
  adrs_buf( 708) <= x"000195c";
  adrs_buf( 709) <= x"000195e";
  adrs_buf( 710) <= x"0001960";
  adrs_buf( 711) <= x"0001962";
  adrs_buf( 712) <= x"0001964";
  adrs_buf( 713) <= x"0001966";
  adrs_buf( 714) <= x"0001968";
  adrs_buf( 715) <= x"000196a";
  adrs_buf( 716) <= x"000196c";
  adrs_buf( 717) <= x"000196e";
  adrs_buf( 718) <= x"0001970";
  adrs_buf( 719) <= x"0001972";
  adrs_buf( 720) <= x"0001974";
  adrs_buf( 721) <= x"0001976";
  adrs_buf( 722) <= x"0001978";
  adrs_buf( 723) <= x"000197a";
  adrs_buf( 724) <= x"000197c";
  adrs_buf( 725) <= x"000197e";
  adrs_buf( 726) <= x"0001980";
  adrs_buf( 727) <= x"0001982";
  adrs_buf( 728) <= x"0001984";
  adrs_buf( 729) <= x"0001986";
  adrs_buf( 730) <= x"0001988";
  adrs_buf( 731) <= x"000198a";
  adrs_buf( 732) <= x"000198c";
  adrs_buf( 733) <= x"000198e";
  adrs_buf( 734) <= x"0001990";
  adrs_buf( 735) <= x"0001992";
  adrs_buf( 736) <= x"0001994";
  adrs_buf( 737) <= x"0001996";
  adrs_buf( 738) <= x"0001998";
  adrs_buf( 739) <= x"000199a";
  adrs_buf( 740) <= x"000199c";
  adrs_buf( 741) <= x"000199e";
  adrs_buf( 742) <= x"00019a0";
  adrs_buf( 743) <= x"00019a2";
  adrs_buf( 744) <= x"00019a4";
  adrs_buf( 745) <= x"00019a6";
  adrs_buf( 746) <= x"00019a8";
  adrs_buf( 747) <= x"00019aa";
  adrs_buf( 748) <= x"00019ac";
  adrs_buf( 749) <= x"00019ae";
  adrs_buf( 750) <= x"00019b0";
  adrs_buf( 751) <= x"00019b2";
  adrs_buf( 752) <= x"00019b4";
  adrs_buf( 753) <= x"00019b6";
  adrs_buf( 754) <= x"00019b8";
  adrs_buf( 755) <= x"00019ba";
  adrs_buf( 756) <= x"00019bc";
  adrs_buf( 757) <= x"00019be";
  adrs_buf( 758) <= x"00019c0";
  adrs_buf( 759) <= x"00019c2";
  adrs_buf( 760) <= x"00019c4";
  adrs_buf( 761) <= x"00019c6";
  adrs_buf( 762) <= x"00019c8";
  adrs_buf( 763) <= x"00019ca";
  adrs_buf( 764) <= x"00019cc";
  adrs_buf( 765) <= x"00019ce";
  adrs_buf( 766) <= x"00019d0";
  adrs_buf( 767) <= x"00019d2";
  adrs_buf( 768) <= x"00019d4";
  adrs_buf( 769) <= x"00019d6";
  adrs_buf( 770) <= x"00019d8";
  adrs_buf( 771) <= x"00019da";
  adrs_buf( 772) <= x"00019dc";
  adrs_buf( 773) <= x"00019de";
  adrs_buf( 774) <= x"00019e0";
  adrs_buf( 775) <= x"00019e2";
  adrs_buf( 776) <= x"00019e4";
  adrs_buf( 777) <= x"00019e6";
  adrs_buf( 778) <= x"00019e8";
  adrs_buf( 779) <= x"00019ea";
  adrs_buf( 780) <= x"00019ec";
  adrs_buf( 781) <= x"00019ee";
  adrs_buf( 782) <= x"00019f0";
  adrs_buf( 783) <= x"00019f2";
  adrs_buf( 784) <= x"00019f4";
  adrs_buf( 785) <= x"00019f6";
  adrs_buf( 786) <= x"00019f8";
  adrs_buf( 787) <= x"00019fa";
  adrs_buf( 788) <= x"00019fc";
  adrs_buf( 789) <= x"00019fe";
  adrs_buf( 790) <= x"0001a00";
  adrs_buf( 791) <= x"0001a02";
  adrs_buf( 792) <= x"0001a04";
  adrs_buf( 793) <= x"0001a06";
  adrs_buf( 794) <= x"0001a08";
  adrs_buf( 795) <= x"0001a0a";
  adrs_buf( 796) <= x"0001a0c";
  adrs_buf( 797) <= x"0001a0e";
  adrs_buf( 798) <= x"0001a10";
  adrs_buf( 799) <= x"0001a12";
  adrs_buf( 800) <= x"0001a14";
  adrs_buf( 801) <= x"0001a16";
  adrs_buf( 802) <= x"0001a18";
  adrs_buf( 803) <= x"0001a1a";
  adrs_buf( 804) <= x"0001a1c";
  adrs_buf( 805) <= x"0001a1e";
  adrs_buf( 806) <= x"0001a20";
  adrs_buf( 807) <= x"0001a22";
  adrs_buf( 808) <= x"0001a24";
  adrs_buf( 809) <= x"0001a26";
  adrs_buf( 810) <= x"0001a28";
  adrs_buf( 811) <= x"0001a2a";
  adrs_buf( 812) <= x"0001a2c";
  adrs_buf( 813) <= x"0001a2e";
  adrs_buf( 814) <= x"0001a30";
  adrs_buf( 815) <= x"0001a32";
  adrs_buf( 816) <= x"0001a34";
  adrs_buf( 817) <= x"0001a36";
  adrs_buf( 818) <= x"0001a38";
  adrs_buf( 819) <= x"0001a3a";
  adrs_buf( 820) <= x"0001a3c";
  adrs_buf( 821) <= x"0001a3e";
  adrs_buf( 822) <= x"0001a40";
  adrs_buf( 823) <= x"0001a42";
  adrs_buf( 824) <= x"0001a44";
  adrs_buf( 825) <= x"0001a46";
  adrs_buf( 826) <= x"0001a48";
  adrs_buf( 827) <= x"0001a4a";
  adrs_buf( 828) <= x"0001a4c";
  adrs_buf( 829) <= x"0001a4e";
  adrs_buf( 830) <= x"0001a50";
  adrs_buf( 831) <= x"0001a52";
  adrs_buf( 832) <= x"0001a54";
  adrs_buf( 833) <= x"0001a56";
  adrs_buf( 834) <= x"0001a58";
  adrs_buf( 835) <= x"0001a5a";
  adrs_buf( 836) <= x"0001a5c";
  adrs_buf( 837) <= x"0001a5e";
  adrs_buf( 838) <= x"0001a60";
  adrs_buf( 839) <= x"0001a62";
  adrs_buf( 840) <= x"0001a64";
  adrs_buf( 841) <= x"0001a66";
  adrs_buf( 842) <= x"0001a68";
  adrs_buf( 843) <= x"0001a6a";
  adrs_buf( 844) <= x"0001a6c";
  adrs_buf( 845) <= x"0001a6e";
  adrs_buf( 846) <= x"0001a70";
  adrs_buf( 847) <= x"0001a72";
  adrs_buf( 848) <= x"0001a74";
  adrs_buf( 849) <= x"0001a76";
  adrs_buf( 850) <= x"0001a78";
  adrs_buf( 851) <= x"0001a7a";
  adrs_buf( 852) <= x"0001a7c";
  adrs_buf( 853) <= x"0001a7e";
  adrs_buf( 854) <= x"0001a80";
  adrs_buf( 855) <= x"0001a82";
  adrs_buf( 856) <= x"0001a84";
  adrs_buf( 857) <= x"0001a86";
  adrs_buf( 858) <= x"0001a88";
  adrs_buf( 859) <= x"0001a8a";
  adrs_buf( 860) <= x"0001a8c";
  adrs_buf( 861) <= x"0001a8e";
  adrs_buf( 862) <= x"0001a90";
  adrs_buf( 863) <= x"0001a92";
  adrs_buf( 864) <= x"0001a94";
  adrs_buf( 865) <= x"0001a96";
  adrs_buf( 866) <= x"0001a98";
  adrs_buf( 867) <= x"0001a9a";
  adrs_buf( 868) <= x"0001a9c";
  adrs_buf( 869) <= x"0001a9e";
  adrs_buf( 870) <= x"0001aa0";
  adrs_buf( 871) <= x"0001aa2";
  adrs_buf( 872) <= x"0001aa4";
  adrs_buf( 873) <= x"0001aa6";
  adrs_buf( 874) <= x"0001aa8";
  adrs_buf( 875) <= x"0001aaa";
  adrs_buf( 876) <= x"0001aac";
  adrs_buf( 877) <= x"0001aae";
  adrs_buf( 878) <= x"0001ab0";
  adrs_buf( 879) <= x"0001ab2";
  adrs_buf( 880) <= x"0001ab4";
  adrs_buf( 881) <= x"0001ab6";
  adrs_buf( 882) <= x"0001ab8";
  adrs_buf( 883) <= x"0001aba";
  adrs_buf( 884) <= x"0001abc";
  adrs_buf( 885) <= x"0001abe";
  adrs_buf( 886) <= x"0001ac0";
  adrs_buf( 887) <= x"0001ac2";
  adrs_buf( 888) <= x"0001ac4";
  adrs_buf( 889) <= x"0001ac6";
  adrs_buf( 890) <= x"0001ac8";
  adrs_buf( 891) <= x"0001aca";
  adrs_buf( 892) <= x"0001acc";
  adrs_buf( 893) <= x"0001ace";
  adrs_buf( 894) <= x"0001ad0";
  adrs_buf( 895) <= x"0001ad2";
  adrs_buf( 896) <= x"0001ad4";
  adrs_buf( 897) <= x"0001ad6";
  adrs_buf( 898) <= x"0001ad8";
  adrs_buf( 899) <= x"0001ada";
  adrs_buf( 900) <= x"0001adc";
  adrs_buf( 901) <= x"0001ade";
  adrs_buf( 902) <= x"0001ae0";
  adrs_buf( 903) <= x"0001ae2";
  adrs_buf( 904) <= x"0001ae4";
  adrs_buf( 905) <= x"0001ae6";
  adrs_buf( 906) <= x"0001ae8";
  adrs_buf( 907) <= x"0001aea";
  adrs_buf( 908) <= x"0001aec";
  adrs_buf( 909) <= x"0001aee";
  adrs_buf( 910) <= x"0001af0";
  adrs_buf( 911) <= x"0001af2";
  adrs_buf( 912) <= x"0001af4";
  adrs_buf( 913) <= x"0001af6";
  adrs_buf( 914) <= x"0001af8";
  adrs_buf( 915) <= x"0001afa";
  adrs_buf( 916) <= x"0001afc";
  adrs_buf( 917) <= x"0001afe";
  adrs_buf( 918) <= x"0001b00";
  adrs_buf( 919) <= x"0001b02";
  adrs_buf( 920) <= x"0001b04";
  adrs_buf( 921) <= x"0001b06";
  adrs_buf( 922) <= x"0001b08";
  adrs_buf( 923) <= x"0001b0a";
  adrs_buf( 924) <= x"0001b0c";
  adrs_buf( 925) <= x"0001b0e";
  adrs_buf( 926) <= x"0001b10";
  adrs_buf( 927) <= x"0001b12";
  adrs_buf( 928) <= x"0001b14";
  adrs_buf( 929) <= x"0001b16";
  adrs_buf( 930) <= x"0001b18";
  adrs_buf( 931) <= x"0001b1a";
  adrs_buf( 932) <= x"0001b1c";
  adrs_buf( 933) <= x"0001b1e";
  adrs_buf( 934) <= x"0001b20";
  adrs_buf( 935) <= x"0001b22";
  adrs_buf( 936) <= x"0001b24";
  adrs_buf( 937) <= x"0001b26";
  adrs_buf( 938) <= x"0001b28";
  adrs_buf( 939) <= x"0001b2a";
  adrs_buf( 940) <= x"0001b2c";
  adrs_buf( 941) <= x"0001b2e";
  adrs_buf( 942) <= x"0001b30";
  adrs_buf( 943) <= x"0001b32";
  adrs_buf( 944) <= x"0001b34";
  adrs_buf( 945) <= x"0001b36";
  adrs_buf( 946) <= x"0001b38";
  adrs_buf( 947) <= x"0001b3a";
  adrs_buf( 948) <= x"0001b3c";
  adrs_buf( 949) <= x"0001b3e";
  adrs_buf( 950) <= x"0001b40";
  adrs_buf( 951) <= x"0001b42";
  adrs_buf( 952) <= x"0001b44";
  adrs_buf( 953) <= x"0001b46";
  adrs_buf( 954) <= x"0001b48";
  adrs_buf( 955) <= x"0001b4a";
  adrs_buf( 956) <= x"0001b4c";
  adrs_buf( 957) <= x"0001b4e";
  adrs_buf( 958) <= x"0001b50";
  adrs_buf( 959) <= x"0001b52";
  adrs_buf( 960) <= x"0001b54";
  adrs_buf( 961) <= x"0001b56";
  adrs_buf( 962) <= x"0001b58";
  adrs_buf( 963) <= x"0001b5a";
  adrs_buf( 964) <= x"0001bb0";
  adrs_buf( 965) <= x"0001bb2";
  adrs_buf( 966) <= x"0001bb4";
  adrs_buf( 967) <= x"0001bb6";
  adrs_buf( 968) <= x"0001bb8";
  adrs_buf( 969) <= x"0001bba";
  adrs_buf( 970) <= x"0000132";
  adrs_buf( 971) <= x"0000134";
  adrs_buf( 972) <= x"0000136";
  adrs_buf( 973) <= x"0001be0";
  adrs_buf( 974) <= x"0001be2";
  adrs_buf( 975) <= x"0001be4";
  adrs_buf( 976) <= x"0001bf4";
  adrs_buf( 977) <= x"0001bf6";
  adrs_buf( 978) <= x"0001bf8";
  adrs_buf( 979) <= x"0001bfa";
  adrs_buf( 980) <= x"0001bfc";
  adrs_buf( 981) <= x"0001bfe";
  adrs_buf( 982) <= x"0001c00";
  adrs_buf( 983) <= x"0001c02";
  adrs_buf( 984) <= x"0001c04";
  adrs_buf( 985) <= x"0001c06";
  adrs_buf( 986) <= x"0001c08";
  adrs_buf( 987) <= x"0001c0a";
  adrs_buf( 988) <= x"0001c0c";
  adrs_buf( 989) <= x"0001c0e";
  adrs_buf( 990) <= x"0001c10";
  adrs_buf( 991) <= x"0001c12";
  adrs_buf( 992) <= x"0001c14";
  adrs_buf( 993) <= x"0001c16";
  adrs_buf( 994) <= x"0001c18";
  adrs_buf( 995) <= x"0001c1a";
  adrs_buf( 996) <= x"0001c1c";
  adrs_buf( 997) <= x"0001c1e";
  adrs_buf( 998) <= x"0001c20";
  adrs_buf( 999) <= x"0001c22";
  --
  adrs_buf(1000) <= x"0001c24";
  adrs_buf(1001) <= x"0001c26";
  adrs_buf(1002) <= x"0001c28";
  adrs_buf(1003) <= x"0001c2a";
  adrs_buf(1004) <= x"0001c2c";
  adrs_buf(1005) <= x"0001c2e";
  adrs_buf(1006) <= x"0001c30";
  adrs_buf(1007) <= x"0001c32";
  adrs_buf(1008) <= x"0001c34";
  adrs_buf(1009) <= x"0001c36";
  adrs_buf(1010) <= x"0001c38";
  adrs_buf(1011) <= x"0001c3a";
  adrs_buf(1012) <= x"0001c60";
  adrs_buf(1013) <= x"0001c62";
  adrs_buf(1014) <= x"0001c64";
  adrs_buf(1015) <= x"0001c66";
  adrs_buf(1016) <= x"0001c68";
  adrs_buf(1017) <= x"0001c6a";
  adrs_buf(1018) <= x"0001c6c";
  adrs_buf(1019) <= x"0001c6e";
  adrs_buf(1020) <= x"0001c70";
  adrs_buf(1021) <= x"0001c72";
  adrs_buf(1022) <= x"0001c74";
  adrs_buf(1023) <= x"0001c76";
  adrs_buf(1024) <= x"0001c78";
  adrs_buf(1025) <= x"0001c7a";
  adrs_buf(1026) <= x"0001c7c";
  adrs_buf(1027) <= x"0001c7e";
  adrs_buf(1028) <= x"0001c80";
  adrs_buf(1029) <= x"0001c82";
  adrs_buf(1030) <= x"0001c84";
  adrs_buf(1031) <= x"0001c86";
  adrs_buf(1032) <= x"0001c88";
  adrs_buf(1033) <= x"0001c8a";
  adrs_buf(1034) <= x"0001c8c";
  adrs_buf(1035) <= x"0001c8e";
  adrs_buf(1036) <= x"0001c90";
  adrs_buf(1037) <= x"0001c92";
  adrs_buf(1038) <= x"0001c94";
  adrs_buf(1039) <= x"0001c96";
  adrs_buf(1040) <= x"0001c98";
  adrs_buf(1041) <= x"0001c9a";
  adrs_buf(1042) <= x"0001c9c";
  adrs_buf(1043) <= x"0001c9e";
  adrs_buf(1044) <= x"0001ca0";
  adrs_buf(1045) <= x"0001ca2";
  adrs_buf(1046) <= x"0001ca4";
  adrs_buf(1047) <= x"0001ca6";
  adrs_buf(1048) <= x"0001ca8";
  adrs_buf(1049) <= x"0001caa";
  adrs_buf(1050) <= x"0001cac";
  adrs_buf(1051) <= x"0001cae";
  adrs_buf(1052) <= x"0001cb0";
  adrs_buf(1053) <= x"0001cb2";
  adrs_buf(1054) <= x"0001cb4";
  adrs_buf(1055) <= x"0001cb6";
  adrs_buf(1056) <= x"0001cb8";
  adrs_buf(1057) <= x"0001cba";
  adrs_buf(1058) <= x"0001cc4";
  adrs_buf(1059) <= x"0001cc6";
  adrs_buf(1060) <= x"0001cc8";
  adrs_buf(1061) <= x"0001cca";
  adrs_buf(1062) <= x"0001ccc";
  adrs_buf(1063) <= x"0001cce";
  adrs_buf(1064) <= x"0001cd0";
  adrs_buf(1065) <= x"0001cd2";
  adrs_buf(1066) <= x"0001cd4";
  adrs_buf(1067) <= x"0001cd6";
  adrs_buf(1068) <= x"0001cd8";
  adrs_buf(1069) <= x"0001cda";
  adrs_buf(1070) <= x"0001cdc";
  adrs_buf(1071) <= x"0001cde";
  adrs_buf(1072) <= x"0001ce0";
  adrs_buf(1073) <= x"0001ce2";
  adrs_buf(1074) <= x"0001ce4";
  adrs_buf(1075) <= x"0001ce6";
  adrs_buf(1076) <= x"0001ce8";
  adrs_buf(1077) <= x"0001cea";
  adrs_buf(1078) <= x"0001cec";
  adrs_buf(1079) <= x"0001cee";
  adrs_buf(1080) <= x"0001cf0";
  adrs_buf(1081) <= x"0001cf2";
  adrs_buf(1082) <= x"0001cf4";
  adrs_buf(1083) <= x"0001cf6";
  adrs_buf(1084) <= x"0001cf8";
  adrs_buf(1085) <= x"0001cfa";
  adrs_buf(1086) <= x"0001cfc";
  adrs_buf(1087) <= x"0001cfe";
  adrs_buf(1088) <= x"0001d00";
  adrs_buf(1089) <= x"0001d02";
  adrs_buf(1090) <= x"0001d04";
  adrs_buf(1091) <= x"0001d06";
  adrs_buf(1092) <= x"0001d08";
  adrs_buf(1093) <= x"0001d0a";
  adrs_buf(1094) <= x"0001d0c";
  adrs_buf(1095) <= x"0001d0e";
  adrs_buf(1096) <= x"0001d10";
  adrs_buf(1097) <= x"0001d12";
  adrs_buf(1098) <= x"0001d14";
  adrs_buf(1099) <= x"0001d16";
  adrs_buf(1100) <= x"0001d18";
  adrs_buf(1101) <= x"0001d1a";
  adrs_buf(1102) <= x"0001d1c";
  adrs_buf(1103) <= x"0001d1e";
  adrs_buf(1104) <= x"0001d20";
  adrs_buf(1105) <= x"0001d22";
  adrs_buf(1106) <= x"0001d24";
  adrs_buf(1107) <= x"0001d1c";
  adrs_buf(1108) <= x"0001d1e";
  adrs_buf(1109) <= x"0001d20";
  adrs_buf(1110) <= x"0001d22";
  adrs_buf(1111) <= x"0001d24";
  adrs_buf(1112) <= x"0001d1c";
  adrs_buf(1113) <= x"0001d1e";
  adrs_buf(1114) <= x"0001d20";
  adrs_buf(1115) <= x"0001d22";
  adrs_buf(1116) <= x"0001d24";
  adrs_buf(1117) <= x"0001d1c";
  adrs_buf(1118) <= x"0001d1e";
  adrs_buf(1119) <= x"0001d20";
  adrs_buf(1120) <= x"0001d22";
  adrs_buf(1121) <= x"0001d24";
  adrs_buf(1122) <= x"0001d1c";
  adrs_buf(1123) <= x"0001d1e";
  adrs_buf(1124) <= x"0001d20";
  adrs_buf(1125) <= x"0001d22";
  adrs_buf(1126) <= x"0001d24";
  adrs_buf(1127) <= x"0001d1c";
  adrs_buf(1128) <= x"0001d1e";
  adrs_buf(1129) <= x"0001d20";
  adrs_buf(1130) <= x"0001d22";
  adrs_buf(1131) <= x"0001d24";
  adrs_buf(1132) <= x"0001d1c";
  adrs_buf(1133) <= x"0001d1e";
  adrs_buf(1134) <= x"0001d20";
  adrs_buf(1135) <= x"0001d22";
  adrs_buf(1136) <= x"0001d24";
  adrs_buf(1137) <= x"0001d1c";
  adrs_buf(1138) <= x"0001d1e";
  adrs_buf(1139) <= x"0001d20";
  adrs_buf(1140) <= x"0001d22";
  adrs_buf(1141) <= x"0001d24";
  adrs_buf(1142) <= x"0001d1c";
  adrs_buf(1143) <= x"0001d1e";
  adrs_buf(1144) <= x"0001d20";
  adrs_buf(1145) <= x"0001d22";
  adrs_buf(1146) <= x"0001d24";
  adrs_buf(1147) <= x"0001d1c";
  adrs_buf(1148) <= x"0001d1e";
  adrs_buf(1149) <= x"0001d20";
  adrs_buf(1150) <= x"0001d22";
  adrs_buf(1151) <= x"0001d24";
  adrs_buf(1152) <= x"0001d26";
  adrs_buf(1153) <= x"0001d28";
  adrs_buf(1154) <= x"0001d2a";
  adrs_buf(1155) <= x"0001d2c";
  adrs_buf(1156) <= x"0001d2e";
  adrs_buf(1157) <= x"0001d30";
  adrs_buf(1158) <= x"0001d32";
  adrs_buf(1159) <= x"0001d34";
  adrs_buf(1160) <= x"0001d36";
  adrs_buf(1161) <= x"0001d38";
  adrs_buf(1162) <= x"0001d3a";
  adrs_buf(1163) <= x"0001d3c";
  adrs_buf(1164) <= x"0001d3e";
  adrs_buf(1165) <= x"0001d40";
  adrs_buf(1166) <= x"0001d42";
  adrs_buf(1167) <= x"0001d44";
  adrs_buf(1168) <= x"0001d46";
  adrs_buf(1169) <= x"0001d48";
  adrs_buf(1170) <= x"0001d4a";
  adrs_buf(1171) <= x"0001d4c";
  adrs_buf(1172) <= x"0001d4e";
  adrs_buf(1173) <= x"0001d50";
  adrs_buf(1174) <= x"0001d52";
  adrs_buf(1175) <= x"0001d54";
  adrs_buf(1176) <= x"0001d56";
  adrs_buf(1177) <= x"0001d58";
  adrs_buf(1178) <= x"0001d5a";
  adrs_buf(1179) <= x"0001d5c";
  adrs_buf(1180) <= x"0001d5e";
  adrs_buf(1181) <= x"0001d60";
  adrs_buf(1182) <= x"0001d62";
  adrs_buf(1183) <= x"0001d64";
  adrs_buf(1184) <= x"0001d66";
  adrs_buf(1185) <= x"0001d68";
  adrs_buf(1186) <= x"0001d6a";
  adrs_buf(1187) <= x"0001d6c";
  adrs_buf(1188) <= x"0001d6e";
  adrs_buf(1189) <= x"0001d70";
  adrs_buf(1190) <= x"0001d72";
  adrs_buf(1191) <= x"0001d74";
  adrs_buf(1192) <= x"0001d76";
  adrs_buf(1193) <= x"0001d78";
  adrs_buf(1194) <= x"0001d7a";
  adrs_buf(1195) <= x"0001d7c";
  adrs_buf(1196) <= x"0001d7e";
  adrs_buf(1197) <= x"0001d80";
  adrs_buf(1198) <= x"0001d82";
  adrs_buf(1199) <= x"0001d84";
  adrs_buf(1200) <= x"0001d86";
  adrs_buf(1201) <= x"0001d88";
  adrs_buf(1202) <= x"0001d8a";
  adrs_buf(1203) <= x"0001d8c";
  adrs_buf(1204) <= x"0001d8e";
  adrs_buf(1205) <= x"0001d90";
  adrs_buf(1206) <= x"0001d92";
  adrs_buf(1207) <= x"0001d94";
  adrs_buf(1208) <= x"0001d96";
  adrs_buf(1209) <= x"0001d98";
  adrs_buf(1210) <= x"0001d9a";
  adrs_buf(1211) <= x"0001d9c";
  adrs_buf(1212) <= x"0001d9e";
  adrs_buf(1213) <= x"0001da0";
  adrs_buf(1214) <= x"0001da2";
  adrs_buf(1215) <= x"0001da4";
  adrs_buf(1216) <= x"0001da6";
  adrs_buf(1217) <= x"0001da8";
  adrs_buf(1218) <= x"0001daa";
  adrs_buf(1219) <= x"0001dac";
  adrs_buf(1220) <= x"0001dae";
  adrs_buf(1221) <= x"0001db0";
  adrs_buf(1222) <= x"0001db2";
  adrs_buf(1223) <= x"0001db4";
  adrs_buf(1224) <= x"0001db6";
  adrs_buf(1225) <= x"0001db8";
  adrs_buf(1226) <= x"0001dba";
  adrs_buf(1227) <= x"0001dbc";
  adrs_buf(1228) <= x"0001dbe";
  adrs_buf(1229) <= x"0001dc0";
  adrs_buf(1230) <= x"0001dc2";
  adrs_buf(1231) <= x"0001dc4";
  adrs_buf(1232) <= x"0001dc6";
  adrs_buf(1233) <= x"0001dc8";
  adrs_buf(1234) <= x"0001dca";
  adrs_buf(1235) <= x"0001dcc";
  adrs_buf(1236) <= x"0001dce";
  adrs_buf(1237) <= x"0001dd0";
  adrs_buf(1238) <= x"0001dd2";
  adrs_buf(1239) <= x"0001dd4";
  adrs_buf(1240) <= x"0001dd6";
  adrs_buf(1241) <= x"0001dd8";
  adrs_buf(1242) <= x"0001dda";
  adrs_buf(1243) <= x"0001ddc";
  adrs_buf(1244) <= x"0001dde";
  adrs_buf(1245) <= x"0001de0";
  adrs_buf(1246) <= x"0001de2";
  adrs_buf(1247) <= x"0001de4";
  adrs_buf(1248) <= x"0001de6";
  adrs_buf(1249) <= x"0001de8";
  adrs_buf(1250) <= x"0001dea";
  adrs_buf(1251) <= x"0001dec";
  adrs_buf(1252) <= x"0001dee";
  adrs_buf(1253) <= x"0001df0";
  adrs_buf(1254) <= x"0001df2";
  adrs_buf(1255) <= x"0001df4";
  adrs_buf(1256) <= x"0001df6";
  adrs_buf(1257) <= x"0001df8";
  adrs_buf(1258) <= x"0001dfa";
  adrs_buf(1259) <= x"0001dfc";
  adrs_buf(1260) <= x"0001dfe";
  adrs_buf(1261) <= x"0001e00";
  adrs_buf(1262) <= x"0001e02";
  adrs_buf(1263) <= x"0001e04";
  adrs_buf(1264) <= x"0001e06";
  adrs_buf(1265) <= x"0001e08";
  adrs_buf(1266) <= x"0001e0a";
  adrs_buf(1267) <= x"0001e0c";
  adrs_buf(1268) <= x"0001e0e";
  adrs_buf(1269) <= x"0001e10";
  adrs_buf(1270) <= x"0001e12";
  adrs_buf(1271) <= x"0001e14";
  adrs_buf(1272) <= x"0001e16";
  adrs_buf(1273) <= x"0001e18";
  adrs_buf(1274) <= x"0001e1a";
  adrs_buf(1275) <= x"0001e1c";
  adrs_buf(1276) <= x"0001e1e";
  adrs_buf(1277) <= x"0001e20";
  adrs_buf(1278) <= x"0001e22";
  adrs_buf(1279) <= x"0001e24";
  adrs_buf(1280) <= x"0001e26";
  adrs_buf(1281) <= x"0001e28";
  adrs_buf(1282) <= x"0001e2a";
  adrs_buf(1283) <= x"0001e2c";
  adrs_buf(1284) <= x"0001e2e";
  adrs_buf(1285) <= x"0001e30";
  adrs_buf(1286) <= x"0001e32";
  adrs_buf(1287) <= x"0001e34";
  adrs_buf(1288) <= x"0001e36";
  adrs_buf(1289) <= x"0001e38";
  adrs_buf(1290) <= x"0001e3a";
  adrs_buf(1291) <= x"0001e3c";
  adrs_buf(1292) <= x"0001e3e";
  adrs_buf(1293) <= x"0001e40";
  adrs_buf(1294) <= x"0001e42";
  adrs_buf(1295) <= x"0001e44";
  adrs_buf(1296) <= x"0001e46";
  adrs_buf(1297) <= x"0001e48";
  adrs_buf(1298) <= x"0001e4a";
  adrs_buf(1299) <= x"0001e4c";
  adrs_buf(1300) <= x"0001e4e";
  adrs_buf(1301) <= x"0001e50";
  adrs_buf(1302) <= x"0001e52";
  adrs_buf(1303) <= x"0001e54";
  adrs_buf(1304) <= x"0001e56";
  adrs_buf(1305) <= x"0001e58";
  adrs_buf(1306) <= x"0001e5a";
  adrs_buf(1307) <= x"0001e5c";
  adrs_buf(1308) <= x"0001e5e";
  adrs_buf(1309) <= x"0001e60";
  adrs_buf(1310) <= x"0001e62";
  adrs_buf(1311) <= x"0001e64";
  adrs_buf(1312) <= x"0001e66";
  adrs_buf(1313) <= x"0001e68";
  adrs_buf(1314) <= x"0001e6a";
  adrs_buf(1315) <= x"0001e6c";
  adrs_buf(1316) <= x"0001e6e";
  adrs_buf(1317) <= x"0001e70";
  adrs_buf(1318) <= x"0001e72";
  adrs_buf(1319) <= x"0001e74";
  adrs_buf(1320) <= x"0001e76";
  adrs_buf(1321) <= x"0001e78";
  adrs_buf(1322) <= x"0001e7a";
  adrs_buf(1323) <= x"0001e7c";
  adrs_buf(1324) <= x"0001e7e";
  adrs_buf(1325) <= x"0001e80";
  adrs_buf(1326) <= x"0001e82";
  adrs_buf(1327) <= x"0001e84";
  adrs_buf(1328) <= x"0001e86";
  adrs_buf(1329) <= x"0001e88";
  adrs_buf(1330) <= x"0001e8a";
  adrs_buf(1331) <= x"0001e8c";
  adrs_buf(1332) <= x"0001e8e";
  adrs_buf(1333) <= x"0001e90";
  adrs_buf(1334) <= x"0001e92";
  adrs_buf(1335) <= x"0001e94";
  adrs_buf(1336) <= x"0001e96";
  adrs_buf(1337) <= x"0001e98";
  adrs_buf(1338) <= x"0001e9a";
  adrs_buf(1339) <= x"0001e9c";
  adrs_buf(1340) <= x"0001e9e";
  adrs_buf(1341) <= x"0001ea0";
  adrs_buf(1342) <= x"0001ea2";
  adrs_buf(1343) <= x"0001ea4";
  adrs_buf(1344) <= x"0001ea6";
  adrs_buf(1345) <= x"0001ea8";
  adrs_buf(1346) <= x"0001eaa";
  adrs_buf(1347) <= x"0001eac";
  adrs_buf(1348) <= x"0001eae";
  adrs_buf(1349) <= x"0001eb0";
  adrs_buf(1350) <= x"0001eb2";
  adrs_buf(1351) <= x"0001eb4";
  adrs_buf(1352) <= x"0001eb6";
  adrs_buf(1353) <= x"0001eb8";
  adrs_buf(1354) <= x"0001eba";
  adrs_buf(1355) <= x"0001ebc";
  adrs_buf(1356) <= x"0001ebe";
  adrs_buf(1357) <= x"0001ec0";
  adrs_buf(1358) <= x"0001ec2";
  adrs_buf(1359) <= x"0001ec4";
  adrs_buf(1360) <= x"0001ec6";
  adrs_buf(1361) <= x"0001ec8";
  adrs_buf(1362) <= x"0001eca";
  adrs_buf(1363) <= x"0001ecc";
  adrs_buf(1364) <= x"0001ece";
  adrs_buf(1365) <= x"0001ed0";
  adrs_buf(1366) <= x"0001ed2";
  adrs_buf(1367) <= x"0001ed4";
  adrs_buf(1368) <= x"0001ed6";
  adrs_buf(1369) <= x"0001ed8";
  adrs_buf(1370) <= x"0001eda";
  adrs_buf(1371) <= x"0001edc";
  adrs_buf(1372) <= x"0001ede";
  adrs_buf(1373) <= x"0001ee0";
  adrs_buf(1374) <= x"0001ee2";
  adrs_buf(1375) <= x"0001ee4";
  adrs_buf(1376) <= x"0001ee6";
  adrs_buf(1377) <= x"0001ee8";
  adrs_buf(1378) <= x"0001eea";
  adrs_buf(1379) <= x"0001eec";
  adrs_buf(1380) <= x"0001eee";
  adrs_buf(1381) <= x"0001ef0";
  adrs_buf(1382) <= x"0001ef2";
  adrs_buf(1383) <= x"0001ef4";
  adrs_buf(1384) <= x"0001ef6";
  adrs_buf(1385) <= x"0001ef8";
  adrs_buf(1386) <= x"0001efa";
  adrs_buf(1387) <= x"0001efc";
  adrs_buf(1388) <= x"0001efe";
  adrs_buf(1389) <= x"0001f00";
  adrs_buf(1390) <= x"0001f02";
  adrs_buf(1391) <= x"0001f04";
  adrs_buf(1392) <= x"0001f06";
  adrs_buf(1393) <= x"0001f08";
  adrs_buf(1394) <= x"0001f0a";
  adrs_buf(1395) <= x"0001f0c";
  adrs_buf(1396) <= x"0001f0e";
  adrs_buf(1397) <= x"0001f10";
  adrs_buf(1398) <= x"0001f12";
  adrs_buf(1399) <= x"0001f14";
  adrs_buf(1400) <= x"0001f16";
  adrs_buf(1401) <= x"0001f18";
  adrs_buf(1402) <= x"0001f1a";
  adrs_buf(1403) <= x"0001f1c";
  adrs_buf(1404) <= x"0001f1e";
  adrs_buf(1405) <= x"0001f20";
  adrs_buf(1406) <= x"0001f22";
  adrs_buf(1407) <= x"0001f24";
  adrs_buf(1408) <= x"0001f26";
  adrs_buf(1409) <= x"0001f28";
  adrs_buf(1410) <= x"0001f2a";
  adrs_buf(1411) <= x"0001f2c";
  adrs_buf(1412) <= x"0001f2e";
  adrs_buf(1413) <= x"0001f30";
  adrs_buf(1414) <= x"0001f32";
  adrs_buf(1415) <= x"0001f34";
  adrs_buf(1416) <= x"0001f36";
  adrs_buf(1417) <= x"0001f38";
  adrs_buf(1418) <= x"0001f3a";
  adrs_buf(1419) <= x"0001f3c";
  adrs_buf(1420) <= x"0001f3e";
  adrs_buf(1421) <= x"0001f40";
  adrs_buf(1422) <= x"0001f42";
  adrs_buf(1423) <= x"0001f44";
  adrs_buf(1424) <= x"0001f46";
  adrs_buf(1425) <= x"0001f48";
  adrs_buf(1426) <= x"0001f4a";
  adrs_buf(1427) <= x"0001f4c";
  adrs_buf(1428) <= x"0001f4e";
  adrs_buf(1429) <= x"0001f50";
  adrs_buf(1430) <= x"0001f52";
  adrs_buf(1431) <= x"0001f54";
  adrs_buf(1432) <= x"0001f56";
  adrs_buf(1433) <= x"0001f58";
  adrs_buf(1434) <= x"0001f5a";
  adrs_buf(1435) <= x"0001f5c";
  adrs_buf(1436) <= x"0001f5e";
  adrs_buf(1437) <= x"0001f60";
  adrs_buf(1438) <= x"0001f62";
  adrs_buf(1439) <= x"0001f64";
  adrs_buf(1440) <= x"0001f66";
  adrs_buf(1441) <= x"0001f68";
  adrs_buf(1442) <= x"0001f6a";
  adrs_buf(1443) <= x"0001f6c";
  adrs_buf(1444) <= x"0001f6e";
  adrs_buf(1445) <= x"0001f70";
  adrs_buf(1446) <= x"0001f72";
  adrs_buf(1447) <= x"0001f74";
  adrs_buf(1448) <= x"0001f76";
  adrs_buf(1449) <= x"0001f78";
  adrs_buf(1450) <= x"0001f7a";
  adrs_buf(1451) <= x"0001f7c";
  adrs_buf(1452) <= x"0001f7e";
  adrs_buf(1453) <= x"0001f80";
  adrs_buf(1454) <= x"0001f82";
  adrs_buf(1455) <= x"0001f84";
  adrs_buf(1456) <= x"0001f86";
  adrs_buf(1457) <= x"0001f88";
  adrs_buf(1458) <= x"0001f8a";
  adrs_buf(1459) <= x"0001f8c";
  adrs_buf(1460) <= x"0001f8e";
  adrs_buf(1461) <= x"0001f90";
  adrs_buf(1462) <= x"0001f92";
  adrs_buf(1463) <= x"0001f94";
  adrs_buf(1464) <= x"0001f96";
  adrs_buf(1465) <= x"0001f98";
  adrs_buf(1466) <= x"0001f9a";
  adrs_buf(1467) <= x"0001f9c";
  adrs_buf(1468) <= x"0001f9e";
  adrs_buf(1469) <= x"0001fa0";
  adrs_buf(1470) <= x"0001fa2";
  adrs_buf(1471) <= x"0001fa4";
  adrs_buf(1472) <= x"0001fa6";
  adrs_buf(1473) <= x"0001fa8";
  adrs_buf(1474) <= x"0001faa";
  adrs_buf(1475) <= x"0001fac";
  adrs_buf(1476) <= x"0001fae";
  adrs_buf(1477) <= x"0001fb0";
  adrs_buf(1478) <= x"0001fb2";
  adrs_buf(1479) <= x"0001fb4";
  adrs_buf(1480) <= x"0001fb6";
  adrs_buf(1481) <= x"0001fb8";
  adrs_buf(1482) <= x"0001fba";
  adrs_buf(1483) <= x"0001fbc";
  adrs_buf(1484) <= x"0001fbe";
  adrs_buf(1485) <= x"0001fc0";
  adrs_buf(1486) <= x"0001fc2";
  adrs_buf(1487) <= x"0001fc4";
  adrs_buf(1488) <= x"0001fc6";
  adrs_buf(1489) <= x"0001fc8";
  adrs_buf(1490) <= x"0001fca";
  adrs_buf(1491) <= x"0001fcc";
  adrs_buf(1492) <= x"0001fce";
  adrs_buf(1493) <= x"0001fd0";
  adrs_buf(1494) <= x"0001fd2";
  adrs_buf(1495) <= x"0001fd4";
  adrs_buf(1496) <= x"0001fd6";
  adrs_buf(1497) <= x"0001fd8";
  adrs_buf(1498) <= x"0001fda";
  adrs_buf(1499) <= x"0001fdc";
  adrs_buf(1500) <= x"0001fde";
  adrs_buf(1501) <= x"0001fe0";
  adrs_buf(1502) <= x"0001fe2";
  adrs_buf(1503) <= x"0001fe4";
  adrs_buf(1504) <= x"0001fe6";
  adrs_buf(1505) <= x"0001fe8";
  adrs_buf(1506) <= x"0001fea";
  adrs_buf(1507) <= x"0001fec";
  adrs_buf(1508) <= x"0001fee";
  adrs_buf(1509) <= x"0001ff0";
  adrs_buf(1510) <= x"0001ff2";
  adrs_buf(1511) <= x"0001ff4";
  adrs_buf(1512) <= x"0001ff6";
  adrs_buf(1513) <= x"0001ff8";
  adrs_buf(1514) <= x"0001ffa";
  adrs_buf(1515) <= x"0001ffc";
  adrs_buf(1516) <= x"0001ffe";
  adrs_buf(1517) <= x"0002000";
  adrs_buf(1518) <= x"0002002";
  adrs_buf(1519) <= x"0002004";
  adrs_buf(1520) <= x"0002006";
  adrs_buf(1521) <= x"0002008";
  adrs_buf(1522) <= x"000200a";
  adrs_buf(1523) <= x"000200c";
  adrs_buf(1524) <= x"000200e";
  adrs_buf(1525) <= x"0002010";
  adrs_buf(1526) <= x"0002012";
  adrs_buf(1527) <= x"0002014";
  adrs_buf(1528) <= x"0002016";
  adrs_buf(1529) <= x"0002018";
  adrs_buf(1530) <= x"000201a";
  adrs_buf(1531) <= x"000201c";
  adrs_buf(1532) <= x"000201e";
  adrs_buf(1533) <= x"0002020";
  adrs_buf(1534) <= x"0002022";
  adrs_buf(1535) <= x"0002024";
  adrs_buf(1536) <= x"0002026";
  adrs_buf(1537) <= x"0002028";
  adrs_buf(1538) <= x"000202a";
  adrs_buf(1539) <= x"000202c";
  adrs_buf(1540) <= x"000202e";
  adrs_buf(1541) <= x"0002030";
  adrs_buf(1542) <= x"0002064";
  adrs_buf(1543) <= x"0002066";
  adrs_buf(1544) <= x"0002068";
  adrs_buf(1545) <= x"000206a";
  adrs_buf(1546) <= x"000206c";
  adrs_buf(1547) <= x"0000138";
  adrs_buf(1548) <= x"000013a";
  adrs_buf(1549) <= x"000013c";
  adrs_buf(1550) <= x"0002090";
  adrs_buf(1551) <= x"0002092";
  adrs_buf(1552) <= x"0002094";
  adrs_buf(1553) <= x"0002096";
  adrs_buf(1554) <= x"000209c";
  adrs_buf(1555) <= x"000209e";
  adrs_buf(1556) <= x"00020a0";
  adrs_buf(1557) <= x"00020a2";
  adrs_buf(1558) <= x"00020a4";
  adrs_buf(1559) <= x"00020a6";
  adrs_buf(1560) <= x"00020a8";
  adrs_buf(1561) <= x"00020aa";
  adrs_buf(1562) <= x"00020ac";
  adrs_buf(1563) <= x"00020ae";
  adrs_buf(1564) <= x"00020b0";
  adrs_buf(1565) <= x"00020b2";
  adrs_buf(1566) <= x"00020b4";
  adrs_buf(1567) <= x"00020b6";
  adrs_buf(1568) <= x"00020b8";
  adrs_buf(1569) <= x"00020ba";
  adrs_buf(1570) <= x"00020bc";
  adrs_buf(1571) <= x"00020be";
  adrs_buf(1572) <= x"00020c0";
  adrs_buf(1573) <= x"00020c2";
  adrs_buf(1574) <= x"00020c4";
  adrs_buf(1575) <= x"00020c6";
  adrs_buf(1576) <= x"00020c8";
  adrs_buf(1577) <= x"00020ca";
  adrs_buf(1578) <= x"00020cc";
  adrs_buf(1579) <= x"00020ce";
  adrs_buf(1580) <= x"00020d0";
  adrs_buf(1581) <= x"00020d2";
  adrs_buf(1582) <= x"00020d4";
  adrs_buf(1583) <= x"00020d6";
  adrs_buf(1584) <= x"00020d8";
  adrs_buf(1585) <= x"00020da";
  adrs_buf(1586) <= x"00020dc";
  adrs_buf(1587) <= x"00020de";
  adrs_buf(1588) <= x"00020e0";
  adrs_buf(1589) <= x"00020e2";
  adrs_buf(1590) <= x"00020e4";
  adrs_buf(1591) <= x"00020e6";
  adrs_buf(1592) <= x"00020e8";
  adrs_buf(1593) <= x"00020ea";
  adrs_buf(1594) <= x"00020ec";
  adrs_buf(1595) <= x"00020ee";
  adrs_buf(1596) <= x"00020f0";
  adrs_buf(1597) <= x"00020f2";
  adrs_buf(1598) <= x"00020f4";
  adrs_buf(1599) <= x"00020f6";
  adrs_buf(1600) <= x"00020f8";
  adrs_buf(1601) <= x"00020fa";
  adrs_buf(1602) <= x"00020fc";
  adrs_buf(1603) <= x"00020fe";
  adrs_buf(1604) <= x"0002100";
  adrs_buf(1605) <= x"0002102";
  adrs_buf(1606) <= x"0002104";
  adrs_buf(1607) <= x"0002106";
  adrs_buf(1608) <= x"0002108";
  adrs_buf(1609) <= x"000210a";
  adrs_buf(1610) <= x"000210c";
  adrs_buf(1611) <= x"000210e";
  adrs_buf(1612) <= x"0002110";
  adrs_buf(1613) <= x"0002112";
  adrs_buf(1614) <= x"0002114";
  adrs_buf(1615) <= x"0002116";
  adrs_buf(1616) <= x"0002118";
  adrs_buf(1617) <= x"000211a";
  adrs_buf(1618) <= x"000211c";
  adrs_buf(1619) <= x"000211e";
  adrs_buf(1620) <= x"0002120";
  adrs_buf(1621) <= x"0002122";
  adrs_buf(1622) <= x"0002124";
  adrs_buf(1623) <= x"0002126";
  adrs_buf(1624) <= x"0002128";
  adrs_buf(1625) <= x"000212a";
  adrs_buf(1626) <= x"000212c";
  adrs_buf(1627) <= x"000212e";
  adrs_buf(1628) <= x"0002130";
  adrs_buf(1629) <= x"0002132";
  adrs_buf(1630) <= x"0002134";
  adrs_buf(1631) <= x"0002136";
  adrs_buf(1632) <= x"0002138";
  adrs_buf(1633) <= x"000213a";
  adrs_buf(1634) <= x"000213c";
  adrs_buf(1635) <= x"000213e";
  adrs_buf(1636) <= x"0002140";
  adrs_buf(1637) <= x"0002142";
  adrs_buf(1638) <= x"0002144";
  adrs_buf(1639) <= x"0002146";
  adrs_buf(1640) <= x"0002148";
  adrs_buf(1641) <= x"000214a";
  adrs_buf(1642) <= x"000214c";
  adrs_buf(1643) <= x"000214e";
  adrs_buf(1644) <= x"0002150";
  adrs_buf(1645) <= x"0002152";
  adrs_buf(1646) <= x"0002154";
  adrs_buf(1647) <= x"0002156";
  adrs_buf(1648) <= x"0002158";
  adrs_buf(1649) <= x"000215a";
  adrs_buf(1650) <= x"000215c";
  adrs_buf(1651) <= x"000215e";
  adrs_buf(1652) <= x"0002160";
  adrs_buf(1653) <= x"0002162";
  adrs_buf(1654) <= x"0002164";
  adrs_buf(1655) <= x"0002166";
  adrs_buf(1656) <= x"0002168";
  adrs_buf(1657) <= x"000216a";
  adrs_buf(1658) <= x"000216c";
  adrs_buf(1659) <= x"000216e";
  adrs_buf(1660) <= x"0002170";
  adrs_buf(1661) <= x"0002172";
  adrs_buf(1662) <= x"0002174";
  adrs_buf(1663) <= x"0002176";
  adrs_buf(1664) <= x"0002178";
  adrs_buf(1665) <= x"000217a";
  adrs_buf(1666) <= x"000217c";
  adrs_buf(1667) <= x"000217e";
  adrs_buf(1668) <= x"0002180";
  adrs_buf(1669) <= x"0002182";
  adrs_buf(1670) <= x"0002184";
  adrs_buf(1671) <= x"0002186";
  adrs_buf(1672) <= x"0002188";
  adrs_buf(1673) <= x"000218a";
  adrs_buf(1674) <= x"000218c";
  adrs_buf(1675) <= x"000218e";
  adrs_buf(1676) <= x"0002190";
  adrs_buf(1677) <= x"0002192";
  adrs_buf(1678) <= x"0002194";
  adrs_buf(1679) <= x"0002196";
  adrs_buf(1680) <= x"0002198";
  adrs_buf(1681) <= x"000219a";
  adrs_buf(1682) <= x"000219c";
  adrs_buf(1683) <= x"000219e";
  adrs_buf(1684) <= x"00021a0";
  adrs_buf(1685) <= x"00021a2";
  adrs_buf(1686) <= x"00021a4";
  adrs_buf(1687) <= x"00021a6";
  adrs_buf(1688) <= x"00021a8";
  adrs_buf(1689) <= x"00021aa";
  adrs_buf(1690) <= x"00021ac";
  adrs_buf(1691) <= x"00021ae";
  adrs_buf(1692) <= x"00021b0";
  adrs_buf(1693) <= x"00021b2";
  adrs_buf(1694) <= x"00021b4";
  adrs_buf(1695) <= x"00021b6";
  adrs_buf(1696) <= x"00021b8";
  adrs_buf(1697) <= x"00021ba";
  adrs_buf(1698) <= x"00021bc";
  adrs_buf(1699) <= x"00021be";
  adrs_buf(1700) <= x"00021c0";
  adrs_buf(1701) <= x"00021c2";
  adrs_buf(1702) <= x"00021c4";
  adrs_buf(1703) <= x"00021c6";
  adrs_buf(1704) <= x"00021c8";
  adrs_buf(1705) <= x"00021ca";
  adrs_buf(1706) <= x"00021cc";
  adrs_buf(1707) <= x"00021ce";
  adrs_buf(1708) <= x"00021d0";
  adrs_buf(1709) <= x"00021d2";
  adrs_buf(1710) <= x"00021d4";
  adrs_buf(1711) <= x"00021d6";
  adrs_buf(1712) <= x"00021d8";
  adrs_buf(1713) <= x"00021da";
  adrs_buf(1714) <= x"00021dc";
  adrs_buf(1715) <= x"00021de";
  adrs_buf(1716) <= x"00021e0";
  adrs_buf(1717) <= x"00021e2";
  adrs_buf(1718) <= x"00021e4";
  adrs_buf(1719) <= x"00021e6";
  adrs_buf(1720) <= x"00021e8";
  adrs_buf(1721) <= x"00021ea";
  adrs_buf(1722) <= x"00021ec";
  adrs_buf(1723) <= x"00021ee";
  adrs_buf(1724) <= x"00021f0";
  adrs_buf(1725) <= x"00021f2";
  adrs_buf(1726) <= x"00021f4";
  adrs_buf(1727) <= x"00021f6";
  adrs_buf(1728) <= x"00021f8";
  adrs_buf(1729) <= x"00021fa";
  adrs_buf(1730) <= x"00021fc";
  adrs_buf(1731) <= x"00021fe";
  adrs_buf(1732) <= x"0002200";
  adrs_buf(1733) <= x"0002202";
  adrs_buf(1734) <= x"0002204";
  adrs_buf(1735) <= x"0002206";
  adrs_buf(1736) <= x"0002208";
  adrs_buf(1737) <= x"000220a";
  adrs_buf(1738) <= x"000220c";
  adrs_buf(1739) <= x"000220e";
  adrs_buf(1740) <= x"0002210";
  adrs_buf(1741) <= x"0002212";
  adrs_buf(1742) <= x"0002214";
  adrs_buf(1743) <= x"0002216";
  adrs_buf(1744) <= x"0002218";
  adrs_buf(1745) <= x"000221a";
  adrs_buf(1746) <= x"000221c";
  adrs_buf(1747) <= x"000221e";
  adrs_buf(1748) <= x"0002220";
  adrs_buf(1749) <= x"0002222";
  adrs_buf(1750) <= x"0002224";
  adrs_buf(1751) <= x"0002226";
  adrs_buf(1752) <= x"0002228";
  adrs_buf(1753) <= x"000222a";
  adrs_buf(1754) <= x"000222c";
  adrs_buf(1755) <= x"000222e";
  adrs_buf(1756) <= x"0002230";
  adrs_buf(1757) <= x"0002232";
  adrs_buf(1758) <= x"0002234";
  adrs_buf(1759) <= x"0002236";
  adrs_buf(1760) <= x"0002238";
  adrs_buf(1761) <= x"000223a";
  adrs_buf(1762) <= x"000223c";
  adrs_buf(1763) <= x"000223e";
  adrs_buf(1764) <= x"0002240";
  adrs_buf(1765) <= x"0002242";
  adrs_buf(1766) <= x"0002244";
  adrs_buf(1767) <= x"0002246";
  adrs_buf(1768) <= x"0002248";
  adrs_buf(1769) <= x"000224a";
  adrs_buf(1770) <= x"000224c";
  adrs_buf(1771) <= x"000224e";
  adrs_buf(1772) <= x"0002250";
  adrs_buf(1773) <= x"0002252";
  adrs_buf(1774) <= x"0002254";
  adrs_buf(1775) <= x"0002256";
  adrs_buf(1776) <= x"0002258";
  adrs_buf(1777) <= x"000225a";
  adrs_buf(1778) <= x"000225c";
  adrs_buf(1779) <= x"000225e";
  adrs_buf(1780) <= x"0002260";
  adrs_buf(1781) <= x"0002262";
  adrs_buf(1782) <= x"0002264";
  adrs_buf(1783) <= x"0002266";
  adrs_buf(1784) <= x"0002268";
  adrs_buf(1785) <= x"000226a";
  adrs_buf(1786) <= x"000226c";
  adrs_buf(1787) <= x"000226e";
  adrs_buf(1788) <= x"0002270";
  adrs_buf(1789) <= x"0002272";
  adrs_buf(1790) <= x"0002274";
  adrs_buf(1791) <= x"0002276";
  adrs_buf(1792) <= x"0002278";
  adrs_buf(1793) <= x"000227a";
  adrs_buf(1794) <= x"000227c";
  adrs_buf(1795) <= x"000227e";
  adrs_buf(1796) <= x"0002280";
  adrs_buf(1797) <= x"0002282";
  adrs_buf(1798) <= x"0002284";
  adrs_buf(1799) <= x"0002286";
  adrs_buf(1800) <= x"0002288";
  adrs_buf(1801) <= x"000228a";
  adrs_buf(1802) <= x"000228c";
  adrs_buf(1803) <= x"000228e";
  adrs_buf(1804) <= x"0002290";
  adrs_buf(1805) <= x"0002292";
  adrs_buf(1806) <= x"0002294";
  adrs_buf(1807) <= x"0002296";
  adrs_buf(1808) <= x"0002298";
  adrs_buf(1809) <= x"000229a";
  adrs_buf(1810) <= x"000229c";
  adrs_buf(1811) <= x"000229e";
  adrs_buf(1812) <= x"00022a0";
  adrs_buf(1813) <= x"00022a2";
  adrs_buf(1814) <= x"00022a4";
  adrs_buf(1815) <= x"00022a6";
  adrs_buf(1816) <= x"00022a8";
  adrs_buf(1817) <= x"00022aa";
  adrs_buf(1818) <= x"00022ac";
  adrs_buf(1819) <= x"00022ae";
  adrs_buf(1820) <= x"00022b0";
  adrs_buf(1821) <= x"00022b2";
  adrs_buf(1822) <= x"00022b4";
  adrs_buf(1823) <= x"00022b6";
  adrs_buf(1824) <= x"00022b8";
  adrs_buf(1825) <= x"00022ba";
  adrs_buf(1826) <= x"00022bc";
  adrs_buf(1827) <= x"00022be";
  adrs_buf(1828) <= x"00022c0";
  adrs_buf(1829) <= x"00022c2";
  adrs_buf(1830) <= x"00022c4";
  adrs_buf(1831) <= x"00022c6";
  adrs_buf(1832) <= x"00022c8";
  adrs_buf(1833) <= x"00022ca";
  adrs_buf(1834) <= x"00022cc";
  adrs_buf(1835) <= x"00022ce";
  adrs_buf(1836) <= x"00022d0";
  adrs_buf(1837) <= x"00022d2";
  adrs_buf(1838) <= x"00022d4";
  adrs_buf(1839) <= x"00022d6";
  adrs_buf(1840) <= x"00022d8";
  adrs_buf(1841) <= x"00022da";
  adrs_buf(1842) <= x"00022dc";
  adrs_buf(1843) <= x"00022de";
  adrs_buf(1844) <= x"00022e0";
  adrs_buf(1845) <= x"00022e2";
  adrs_buf(1846) <= x"00022e4";
  adrs_buf(1847) <= x"00022e6";
  adrs_buf(1848) <= x"00022e8";
  adrs_buf(1849) <= x"00022ea";
  adrs_buf(1850) <= x"00022ec";
  adrs_buf(1851) <= x"00022ee";
  adrs_buf(1852) <= x"00022f0";
  adrs_buf(1853) <= x"00022f2";
  adrs_buf(1854) <= x"00022f4";
  adrs_buf(1855) <= x"00022f6";
  adrs_buf(1856) <= x"00022f8";
  adrs_buf(1857) <= x"00022fa";
  adrs_buf(1858) <= x"00022fc";
  adrs_buf(1859) <= x"00022fe";
  adrs_buf(1860) <= x"0002300";
  adrs_buf(1861) <= x"0002302";
  adrs_buf(1862) <= x"0002304";
  adrs_buf(1863) <= x"0002306";
  adrs_buf(1864) <= x"0002308";
  adrs_buf(1865) <= x"000230a";
  adrs_buf(1866) <= x"000230c";
  adrs_buf(1867) <= x"000230e";
  adrs_buf(1868) <= x"0002310";
  adrs_buf(1869) <= x"0002312";
  adrs_buf(1870) <= x"0002314";
  adrs_buf(1871) <= x"0002316";
  adrs_buf(1872) <= x"0002318";
  adrs_buf(1873) <= x"000231a";
  adrs_buf(1874) <= x"000231c";
  adrs_buf(1875) <= x"000231e";
  adrs_buf(1876) <= x"0002320";
  adrs_buf(1877) <= x"0002322";
  adrs_buf(1878) <= x"0002324";
  adrs_buf(1879) <= x"0002326";
  adrs_buf(1880) <= x"0002328";
  adrs_buf(1881) <= x"000232a";
  adrs_buf(1882) <= x"000232c";
  adrs_buf(1883) <= x"000232e";
  adrs_buf(1884) <= x"0002330";
  adrs_buf(1885) <= x"0002332";
  adrs_buf(1886) <= x"0002334";
  adrs_buf(1887) <= x"0002336";
  adrs_buf(1888) <= x"0002338";
  adrs_buf(1889) <= x"000233a";
  adrs_buf(1890) <= x"000233c";
  adrs_buf(1891) <= x"000233e";
  adrs_buf(1892) <= x"0002340";
  adrs_buf(1893) <= x"0002342";
  adrs_buf(1894) <= x"0002344";
  adrs_buf(1895) <= x"0002346";
  adrs_buf(1896) <= x"0002348";
  adrs_buf(1897) <= x"000234a";
  adrs_buf(1898) <= x"000234c";
  adrs_buf(1899) <= x"000234e";
  adrs_buf(1900) <= x"0002350";
  adrs_buf(1901) <= x"0002352";
  adrs_buf(1902) <= x"0002354";
  adrs_buf(1903) <= x"0002356";
  adrs_buf(1904) <= x"0002358";
  adrs_buf(1905) <= x"000235a";
  adrs_buf(1906) <= x"000235c";
  adrs_buf(1907) <= x"000235e";
  adrs_buf(1908) <= x"0002360";
  adrs_buf(1909) <= x"0002362";
  adrs_buf(1910) <= x"0002364";
  adrs_buf(1911) <= x"00024cc";
  adrs_buf(1912) <= x"00024ce";
  adrs_buf(1913) <= x"00024d0";
  adrs_buf(1914) <= x"00024d2";
  adrs_buf(1915) <= x"00024d4";
  adrs_buf(1916) <= x"00024d6";
  adrs_buf(1917) <= x"000013e";
  adrs_buf(1918) <= x"0000140";
  adrs_buf(1919) <= x"0000142";
  adrs_buf(1920) <= x"0002510";
  adrs_buf(1921) <= x"0002512";
  adrs_buf(1922) <= x"0002514";
  adrs_buf(1923) <= x"0002516";
  adrs_buf(1924) <= x"000251c";
  adrs_buf(1925) <= x"000251e";
  adrs_buf(1926) <= x"0002520";
  adrs_buf(1927) <= x"0002522";
  adrs_buf(1928) <= x"0002524";
  adrs_buf(1929) <= x"0002526";
  adrs_buf(1930) <= x"0002528";
  adrs_buf(1931) <= x"000252a";
  adrs_buf(1932) <= x"000252c";
  adrs_buf(1933) <= x"000252e";
  adrs_buf(1934) <= x"0002530";
  adrs_buf(1935) <= x"0002532";
  adrs_buf(1936) <= x"0002534";
  adrs_buf(1937) <= x"0002536";
  adrs_buf(1938) <= x"0002538";
  adrs_buf(1939) <= x"000253a";
  adrs_buf(1940) <= x"000253c";
  adrs_buf(1941) <= x"000253e";
  adrs_buf(1942) <= x"0002540";
  adrs_buf(1943) <= x"0002542";
  adrs_buf(1944) <= x"0002544";
  adrs_buf(1945) <= x"0002546";
  adrs_buf(1946) <= x"0002548";
  adrs_buf(1947) <= x"000254a";
  adrs_buf(1948) <= x"000254c";
  adrs_buf(1949) <= x"000254e";
  adrs_buf(1950) <= x"0002550";
  adrs_buf(1951) <= x"0002552";
  adrs_buf(1952) <= x"0002554";
  adrs_buf(1953) <= x"0002556";
  adrs_buf(1954) <= x"0002558";
  adrs_buf(1955) <= x"000255a";
  adrs_buf(1956) <= x"000255c";
  adrs_buf(1957) <= x"000255e";
  adrs_buf(1958) <= x"0002560";
  adrs_buf(1959) <= x"0002562";
  adrs_buf(1960) <= x"0002564";
  adrs_buf(1961) <= x"0002566";
  adrs_buf(1962) <= x"0002568";
  adrs_buf(1963) <= x"000256a";
  adrs_buf(1964) <= x"000256c";
  adrs_buf(1965) <= x"000256e";
  adrs_buf(1966) <= x"0002570";
  adrs_buf(1967) <= x"00025cc";
  adrs_buf(1968) <= x"00025ce";
  adrs_buf(1969) <= x"00025d0";
  adrs_buf(1970) <= x"00025d2";
  adrs_buf(1971) <= x"00025d4";
  adrs_buf(1972) <= x"00025d6";
  adrs_buf(1973) <= x"00025d8";
  adrs_buf(1974) <= x"00025da";
  adrs_buf(1975) <= x"00025dc";
  adrs_buf(1976) <= x"00025de";
  adrs_buf(1977) <= x"00025e0";
  adrs_buf(1978) <= x"00025e2";
  adrs_buf(1979) <= x"00025e4";
  adrs_buf(1980) <= x"00025e6";
  adrs_buf(1981) <= x"00025e8";
  adrs_buf(1982) <= x"00025ea";
  adrs_buf(1983) <= x"00025ec";
  adrs_buf(1984) <= x"00025ee";
  adrs_buf(1985) <= x"00025f0";
  adrs_buf(1986) <= x"00025f2";
  adrs_buf(1987) <= x"00025f4";
  adrs_buf(1988) <= x"00025f6";
  adrs_buf(1989) <= x"00025f8";
  adrs_buf(1990) <= x"00025fa";
  adrs_buf(1991) <= x"00025fc";
  adrs_buf(1992) <= x"00025fe";
  adrs_buf(1993) <= x"0002600";
  adrs_buf(1994) <= x"0002602";
  adrs_buf(1995) <= x"0002604";
  adrs_buf(1996) <= x"0002606";
  adrs_buf(1997) <= x"0002608";
  adrs_buf(1998) <= x"000260a";
  adrs_buf(1999) <= x"00025dc";
  adrs_buf(2000) <= x"00025de";

end tb;
